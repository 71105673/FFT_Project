`timescale 1ns / 1ps

module tb_fft_top;

    parameter WIDTH = 9;
    parameter WIDTH_DO = 13;

    logic clk, rstn;
    logic fft_mode;
    logic di_en;
    logic signed [WIDTH-1:0] di_re[0:15];
    logic signed [WIDTH-1:0] di_im[0:15];

    logic signed [WIDTH_DO-1:0] do_re[0:15];
    logic signed [WIDTH_DO-1:0] do_im[0:15];

    integer fp;

    // // DUT
    // sdf1 #(
    //     .N(512),
    //     .M(512),
    //     .WIDTH(WIDTH),
    //     .WIDTH_DO(WIDTH_DO)
    // ) dut (
    //     .clk(clk),
    //     .rstn(rstn),
    //     .fft_mode(fft_mode),
    //     .di_en(di_en),
    //     .di_re(di_re),
    //     .di_im(di_im),

    //     .do_index(do_index),
    //     .do_en(do_en),
    //     .do_re(do_re),
    //     .do_im(do_im)
    // );

    fft_top #(
        .WIDTH(9)
    ) dut (
        .clk(clk),
        .rstn(rstn),
        .fft_mode(fft_mode),

        .din_i(di_re),
        .din_q(di_im),
        .din_valid(di_en),

        .do_re(do_re),
        .do_im(do_im),
        .do_en(do_en)
    );

    // Clock
    initial clk = 0;
    always #5 clk = ~clk;

    // Stimulus
    initial begin
        rstn = 0;
        di_en = 0;
        fft_mode = 1;
        #20;
        rstn = 1;
        #10;
        @(posedge clk);
        di_en = 1;
        di_re[0] = 12;
        di_im[0] = 23;
        di_re[1] = 19;
        di_im[1] = 29;
        di_re[2] = 38;
        di_im[2] = 5;
        di_re[3] = 39;
        di_im[3] = 40;
        di_re[4] = 17;
        di_im[4] = 21;
        di_re[5] = 27;
        di_im[5] = 34;
        di_re[6] = 36;
        di_im[6] = 36;
        di_re[7] = 19;
        di_im[7] = 21;
        di_re[8] = 46;
        di_im[8] = 28;
        di_re[9] = 41;
        di_im[9] = 13;
        di_re[10] = 30;
        di_im[10] = 28;
        di_re[11] = 46;
        di_im[11] = 4;
        di_re[12] = 24;
        di_im[12] = 25;
        di_re[13] = 4;
        di_im[13] = 43;
        di_re[14] = 42;
        di_im[14] = 21;
        di_re[15] = 38;
        di_im[15] = 7;

        @(posedge clk);
        di_en = 1;
        di_re[0] = 30;
        di_im[0] = 13;
        di_re[1] = 21;
        di_im[1] = 41;
        di_re[2] = 9;
        di_im[2] = 15;
        di_re[3] = 23;
        di_im[3] = 16;
        di_re[4] = 38;
        di_im[4] = 47;
        di_re[5] = 8;
        di_im[5] = 11;
        di_re[6] = 34;
        di_im[6] = 18;
        di_re[7] = 47;
        di_im[7] = 47;
        di_re[8] = 31;
        di_im[8] = 41;
        di_re[9] = 19;
        di_im[9] = 30;
        di_re[10] = 47;
        di_im[10] = 27;
        di_re[11] = 45;
        di_im[11] = 35;
        di_re[12] = 23;
        di_im[12] = 31;
        di_re[13] = 43;
        di_im[13] = 10;
        di_re[14] = 19;
        di_im[14] = 48;
        di_re[15] = 19;
        di_im[15] = 32;

        @(posedge clk);
        di_en = 1;
        di_re[0] = 43;
        di_im[0] = 48;
        di_re[1] = 31;
        di_im[1] = 5;
        di_re[2] = 2;
        di_im[2] = 30;
        di_re[3] = 27;
        di_im[3] = 46;
        di_re[4] = 36;
        di_im[4] = 32;
        di_re[5] = 25;
        di_im[5] = 12;
        di_re[6] = 46;
        di_im[6] = 26;
        di_re[7] = 1;
        di_im[7] = 33;
        di_re[8] = 25;
        di_im[8] = 3;
        di_re[9] = 43;
        di_im[9] = 16;
        di_re[10] = 11;
        di_im[10] = 5;
        di_re[11] = 15;
        di_im[11] = 11;
        di_re[12] = 31;
        di_im[12] = 3;
        di_re[13] = 13;
        di_im[13] = 14;
        di_re[14] = 42;
        di_im[14] = 21;
        di_re[15] = 36;
        di_im[15] = 29;

        @(posedge clk);
        di_en = 1;
        di_re[0] = 38;
        di_im[0] = 5;
        di_re[1] = 47;
        di_im[1] = 41;
        di_re[2] = 2;
        di_im[2] = 22;
        di_re[3] = 16;
        di_im[3] = 30;
        di_re[4] = 11;
        di_im[4] = 28;
        di_re[5] = 29;
        di_im[5] = 29;
        di_re[6] = 22;
        di_im[6] = 2;
        di_re[7] = 25;
        di_im[7] = 20;
        di_re[8] = 5;
        di_im[8] = 22;
        di_re[9] = 22;
        di_im[9] = 26;
        di_re[10] = 39;
        di_im[10] = 34;
        di_re[11] = 42;
        di_im[11] = 3;
        di_re[12] = 11;
        di_im[12] = 22;
        di_re[13] = 46;
        di_im[13] = 38;
        di_re[14] = 22;
        di_im[14] = 16;
        di_re[15] = 3;
        di_im[15] = 36;

        @(posedge clk);
        di_en = 1;
        di_re[0] = 24;
        di_im[0] = 10;
        di_re[1] = 21;
        di_im[1] = 8;
        di_re[2] = 36;
        di_im[2] = 18;
        di_re[3] = 45;
        di_im[3] = 1;
        di_re[4] = 40;
        di_im[4] = 30;
        di_re[5] = 26;
        di_im[5] = 31;
        di_re[6] = 35;
        di_im[6] = 5;
        di_re[7] = 42;
        di_im[7] = 1;
        di_re[8] = 14;
        di_im[8] = 9;
        di_re[9] = 44;
        di_im[9] = 3;
        di_re[10] = 28;
        di_im[10] = 31;
        di_re[11] = 31;
        di_im[11] = 42;
        di_re[12] = 3;
        di_im[12] = 39;
        di_re[13] = 25;
        di_im[13] = 33;
        di_re[14] = 10;
        di_im[14] = 26;
        di_re[15] = 34;
        di_im[15] = 46;

        @(posedge clk);
        di_en = 1;
        di_re[0] = 21;
        di_im[0] = 4;
        di_re[1] = 3;
        di_im[1] = 30;
        di_re[2] = 38;
        di_im[2] = 33;
        di_re[3] = 17;
        di_im[3] = 45;
        di_re[4] = 25;
        di_im[4] = 46;
        di_re[5] = 4;
        di_im[5] = 10;
        di_re[6] = 37;
        di_im[6] = 44;
        di_re[7] = 38;
        di_im[7] = 14;
        di_re[8] = 7;
        di_im[8] = 41;
        di_re[9] = 38;
        di_im[9] = 13;
        di_re[10] = 11;
        di_im[10] = 15;
        di_re[11] = 40;
        di_im[11] = 39;
        di_re[12] = 27;
        di_im[12] = 27;
        di_re[13] = 14;
        di_im[13] = 34;
        di_re[14] = 38;
        di_im[14] = 21;
        di_re[15] = 21;
        di_im[15] = 22;

        @(posedge clk);
        di_en = 1;
        di_re[0] = 13;
        di_im[0] = 32;
        di_re[1] = 43;
        di_im[1] = 44;
        di_re[2] = 36;
        di_im[2] = 13;
        di_re[3] = 33;
        di_im[3] = 6;
        di_re[4] = 6;
        di_im[4] = 9;
        di_re[5] = 7;
        di_im[5] = 28;
        di_re[6] = 4;
        di_im[6] = 39;
        di_re[7] = 35;
        di_im[7] = 44;
        di_re[8] = 24;
        di_im[8] = 31;
        di_re[9] = 43;
        di_im[9] = 26;
        di_re[10] = 14;
        di_im[10] = 47;
        di_re[11] = 2;
        di_im[11] = 16;
        di_re[12] = 47;
        di_im[12] = 18;
        di_re[13] = 15;
        di_im[13] = 6;
        di_re[14] = 44;
        di_im[14] = 7;
        di_re[15] = 16;
        di_im[15] = 43;

        @(posedge clk);
        di_en = 1;
        di_re[0] = 24;
        di_im[0] = 30;
        di_re[1] = 28;
        di_im[1] = 34;
        di_re[2] = 1;
        di_im[2] = 25;
        di_re[3] = 2;
        di_im[3] = 40;
        di_re[4] = 16;
        di_im[4] = 41;
        di_re[5] = 12;
        di_im[5] = 28;
        di_re[6] = 45;
        di_im[6] = 2;
        di_re[7] = 3;
        di_im[7] = 1;
        di_re[8] = 33;
        di_im[8] = 29;
        di_re[9] = 5;
        di_im[9] = 38;
        di_re[10] = 30;
        di_im[10] = 3;
        di_re[11] = 3;
        di_im[11] = 7;
        di_re[12] = 38;
        di_im[12] = 4;
        di_re[13] = 11;
        di_im[13] = 12;
        di_re[14] = 5;
        di_im[14] = 41;
        di_re[15] = 34;
        di_im[15] = 35;

        @(posedge clk);
        di_en = 1;
        di_re[0] = 31;
        di_im[0] = 25;
        di_re[1] = 16;
        di_im[1] = 32;
        di_re[2] = 6;
        di_im[2] = 7;
        di_re[3] = 1;
        di_im[3] = 46;
        di_re[4] = 47;
        di_im[4] = 6;
        di_re[5] = 22;
        di_im[5] = 32;
        di_re[6] = 14;
        di_im[6] = 36;
        di_re[7] = 27;
        di_im[7] = 21;
        di_re[8] = 13;
        di_im[8] = 36;
        di_re[9] = 43;
        di_im[9] = 35;
        di_re[10] = 20;
        di_im[10] = 45;
        di_re[11] = 12;
        di_im[11] = 26;
        di_re[12] = 46;
        di_im[12] = 13;
        di_re[13] = 12;
        di_im[13] = 45;
        di_re[14] = 3;
        di_im[14] = 14;
        di_re[15] = 28;
        di_im[15] = 10;

        @(posedge clk);
        di_en = 1;
        di_re[0] = 31;
        di_im[0] = 38;
        di_re[1] = 24;
        di_im[1] = 31;
        di_re[2] = 38;
        di_im[2] = 11;
        di_re[3] = 29;
        di_im[3] = 5;
        di_re[4] = 25;
        di_im[4] = 40;
        di_re[5] = 44;
        di_im[5] = 24;
        di_re[6] = 13;
        di_im[6] = 31;
        di_re[7] = 44;
        di_im[7] = 24;
        di_re[8] = 47;
        di_im[8] = 9;
        di_re[9] = 5;
        di_im[9] = 14;
        di_re[10] = 19;
        di_im[10] = 20;
        di_re[11] = 15;
        di_im[11] = 33;
        di_re[12] = 4;
        di_im[12] = 19;
        di_re[13] = 14;
        di_im[13] = 15;
        di_re[14] = 5;
        di_im[14] = 29;
        di_re[15] = 14;
        di_im[15] = 7;

        @(posedge clk);
        di_en = 1;
        di_re[0] = 0;
        di_im[0] = 14;
        di_re[1] = 26;
        di_im[1] = 42;
        di_re[2] = 2;
        di_im[2] = 43;
        di_re[3] = 6;
        di_im[3] = 40;
        di_re[4] = 38;
        di_im[4] = 44;
        di_re[5] = 7;
        di_im[5] = 24;
        di_re[6] = 19;
        di_im[6] = 8;
        di_re[7] = 28;
        di_im[7] = 29;
        di_re[8] = 10;
        di_im[8] = 25;
        di_re[9] = 47;
        di_im[9] = 24;
        di_re[10] = 33;
        di_im[10] = 20;
        di_re[11] = 2;
        di_im[11] = 14;
        di_re[12] = 38;
        di_im[12] = 17;
        di_re[13] = 4;
        di_im[13] = 25;
        di_re[14] = 18;
        di_im[14] = 35;
        di_re[15] = 25;
        di_im[15] = 39;

        @(posedge clk);
        di_en = 1;
        di_re[0] = 39;
        di_im[0] = 9;
        di_re[1] = 6;
        di_im[1] = 39;
        di_re[2] = 31;
        di_im[2] = 1;
        di_re[3] = 43;
        di_im[3] = 25;
        di_re[4] = 26;
        di_im[4] = 29;
        di_re[5] = 37;
        di_im[5] = 41;
        di_re[6] = 18;
        di_im[6] = 4;
        di_re[7] = 35;
        di_im[7] = 16;
        di_re[8] = 40;
        di_im[8] = 18;
        di_re[9] = 40;
        di_im[9] = 8;
        di_re[10] = 6;
        di_im[10] = 42;
        di_re[11] = 2;
        di_im[11] = 33;
        di_re[12] = 35;
        di_im[12] = 21;
        di_re[13] = 18;
        di_im[13] = 47;
        di_re[14] = 19;
        di_im[14] = 21;
        di_re[15] = 8;
        di_im[15] = 16;

        @(posedge clk);
        di_en = 1;
        di_re[0] = 15;
        di_im[0] = 43;
        di_re[1] = 12;
        di_im[1] = 15;
        di_re[2] = 20;
        di_im[2] = 34;
        di_re[3] = 7;
        di_im[3] = 42;
        di_re[4] = 4;
        di_im[4] = 22;
        di_re[5] = 1;
        di_im[5] = 36;
        di_re[6] = 34;
        di_im[6] = 10;
        di_re[7] = 33;
        di_im[7] = 27;
        di_re[8] = 41;
        di_im[8] = 27;
        di_re[9] = 43;
        di_im[9] = 20;
        di_re[10] = 17;
        di_im[10] = 23;
        di_re[11] = 12;
        di_im[11] = 45;
        di_re[12] = 22;
        di_im[12] = 12;
        di_re[13] = 21;
        di_im[13] = 34;
        di_re[14] = 19;
        di_im[14] = 9;
        di_re[15] = 41;
        di_im[15] = 28;

        @(posedge clk);
        di_en = 1;
        di_re[0] = 18;
        di_im[0] = 11;
        di_re[1] = 11;
        di_im[1] = 25;
        di_re[2] = 21;
        di_im[2] = 36;
        di_re[3] = 3;
        di_im[3] = 41;
        di_re[4] = 33;
        di_im[4] = 7;
        di_re[5] = 41;
        di_im[5] = 10;
        di_re[6] = 29;
        di_im[6] = 26;
        di_re[7] = 8;
        di_im[7] = 0;
        di_re[8] = 37;
        di_im[8] = 37;
        di_re[9] = 20;
        di_im[9] = 3;
        di_re[10] = 28;
        di_im[10] = 8;
        di_re[11] = 35;
        di_im[11] = 26;
        di_re[12] = 12;
        di_im[12] = 44;
        di_re[13] = 36;
        di_im[13] = 43;
        di_re[14] = 3;
        di_im[14] = 9;
        di_re[15] = 35;
        di_im[15] = 33;

        @(posedge clk);
        di_en = 1;
        di_re[0] = 37;
        di_im[0] = 24;
        di_re[1] = 20;
        di_im[1] = 29;
        di_re[2] = 41;
        di_im[2] = 32;
        di_re[3] = 25;
        di_im[3] = 14;
        di_re[4] = 34;
        di_im[4] = 18;
        di_re[5] = 27;
        di_im[5] = 43;
        di_re[6] = 40;
        di_im[6] = 43;
        di_re[7] = 45;
        di_im[7] = 39;
        di_re[8] = 0;
        di_im[8] = 0;
        di_re[9] = 4;
        di_im[9] = 13;
        di_re[10] = 1;
        di_im[10] = 20;
        di_re[11] = 16;
        di_im[11] = 26;
        di_re[12] = 44;
        di_im[12] = 14;
        di_re[13] = 16;
        di_im[13] = 41;
        di_re[14] = 16;
        di_im[14] = 7;
        di_re[15] = 24;
        di_im[15] = 41;

        @(posedge clk);
        di_en = 1;
        di_re[0] = 18;
        di_im[0] = 33;
        di_re[1] = 30;
        di_im[1] = 22;
        di_re[2] = 23;
        di_im[2] = 46;
        di_re[3] = 4;
        di_im[3] = 13;
        di_re[4] = 21;
        di_im[4] = 28;
        di_re[5] = 42;
        di_im[5] = 23;
        di_re[6] = 21;
        di_im[6] = 36;
        di_re[7] = 22;
        di_im[7] = 41;
        di_re[8] = 22;
        di_im[8] = 24;
        di_re[9] = 23;
        di_im[9] = 11;
        di_re[10] = 4;
        di_im[10] = 3;
        di_re[11] = 43;
        di_im[11] = 11;
        di_re[12] = 41;
        di_im[12] = 34;
        di_re[13] = 42;
        di_im[13] = 45;
        di_re[14] = 7;
        di_im[14] = 19;
        di_re[15] = 47;
        di_im[15] = 31;

        @(posedge clk);
        di_en = 1;
        di_re[0] = 43;
        di_im[0] = 23;
        di_re[1] = 1;
        di_im[1] = 30;
        di_re[2] = 11;
        di_im[2] = 25;
        di_re[3] = 35;
        di_im[3] = 29;
        di_re[4] = 28;
        di_im[4] = 21;
        di_re[5] = 12;
        di_im[5] = 21;
        di_re[6] = 0;
        di_im[6] = 29;
        di_re[7] = 46;
        di_im[7] = 5;
        di_re[8] = 2;
        di_im[8] = 43;
        di_re[9] = 12;
        di_im[9] = 0;
        di_re[10] = 39;
        di_im[10] = 7;
        di_re[11] = 42;
        di_im[11] = 5;
        di_re[12] = 17;
        di_im[12] = 28;
        di_re[13] = 28;
        di_im[13] = 32;
        di_re[14] = 31;
        di_im[14] = 21;
        di_re[15] = 7;
        di_im[15] = 36;

        @(posedge clk);
        di_en = 1;
        di_re[0] = 12;
        di_im[0] = 31;
        di_re[1] = 41;
        di_im[1] = 4;
        di_re[2] = 47;
        di_im[2] = 2;
        di_re[3] = 40;
        di_im[3] = 40;
        di_re[4] = 2;
        di_im[4] = 26;
        di_re[5] = 45;
        di_im[5] = 15;
        di_re[6] = 39;
        di_im[6] = 29;
        di_re[7] = 38;
        di_im[7] = 38;
        di_re[8] = 2;
        di_im[8] = 14;
        di_re[9] = 31;
        di_im[9] = 24;
        di_re[10] = 47;
        di_im[10] = 36;
        di_re[11] = 27;
        di_im[11] = 14;
        di_re[12] = 12;
        di_im[12] = 43;
        di_re[13] = 21;
        di_im[13] = 39;
        di_re[14] = 5;
        di_im[14] = 41;
        di_re[15] = 1;
        di_im[15] = 43;

	@(posedge clk);
        di_en = 1;
        di_re[0] = 43;
        di_im[0] = 25;
        di_re[1] = 6;
        di_im[1] = 9;
        di_re[2] = 34;
        di_im[2] = 40;
        di_re[3] = 2;
        di_im[3] = 36;
        di_re[4] = 46;
        di_im[4] = 16;
        di_re[5] = 31;
        di_im[5] = 16;
        di_re[6] = 10;
        di_im[6] = 38;
        di_re[7] = 35;
        di_im[7] = 13;
        di_re[8] = 28;
        di_im[8] = 20;
        di_re[9] = 4;
        di_im[9] = 1;
        di_re[10] = 24;
        di_im[10] = 13;
        di_re[11] = 16;
        di_im[11] = 14;
        di_re[12] = 8;
        di_im[12] = 19;
        di_re[13] = 33;
        di_im[13] = 10;
        di_re[14] = 32;
        di_im[14] = 21;
        di_re[15] = 21;
        di_im[15] = 8;

	@(posedge clk);
        di_en = 1;
        di_re[0] = 9;
        di_im[0] = 30;
        di_re[1] = 13;
        di_im[1] = 27;
        di_re[2] = 45;
        di_im[2] = 34;
        di_re[3] = 33;
        di_im[3] = 46;
        di_re[4] = 37;
        di_im[4] = 29;
        di_re[5] = 46;
        di_im[5] = 3;
        di_re[6] = 13;
        di_im[6] = 47;
        di_re[7] = 37;
        di_im[7] = 23;
        di_re[8] = 33;
        di_im[8] = 20;
        di_re[9] = 18;
        di_im[9] = 10;
        di_re[10] = 18;
        di_im[10] = 1;
        di_re[11] = 23;
        di_im[11] = 16;
        di_re[12] = 47;
        di_im[12] = 27;
        di_re[13] = 41;
        di_im[13] = 20;
        di_re[14] = 22;
        di_im[14] = 40;
        di_re[15] = 48;
        di_im[15] = 25;

	@(posedge clk);
	di_en = 1;
        di_re[0] = 44;
        di_im[0] = 35;
        di_re[1] = 27;
        di_im[1] = 47;
        di_re[2] = 40;
        di_im[2] = 46;
        di_re[3] = 31;
        di_im[3] = 18;
        di_re[4] = 23;
        di_im[4] = 44;
        di_re[5] = 1;
        di_im[5] = 8;
        di_re[6] = 23;
        di_im[6] = 26;
        di_re[7] = 3;
        di_im[7] = 32;
        di_re[8] = 43;
        di_im[8] = 5;
        di_re[9] = 21;
        di_im[9] = 13;
        di_re[10] = 47;
        di_im[10] = 29;
        di_re[11] = 12;
        di_im[11] = 6;
        di_re[12] = 26;
        di_im[12] = 40;
        di_re[13] = 40;
        di_im[13] = 40;
        di_re[14] = 10;
        di_im[14] = 26;
        di_re[15] = 42;
        di_im[15] = 6;

        @(posedge clk);
        di_en = 1;
        di_re[0] = 41;
        di_im[0] = 43;
        di_re[1] = 10;
        di_im[1] = 4;
        di_re[2] = 23;
        di_im[2] = 40;
        di_re[3] = 23;
        di_im[3] = 20;
        di_re[4] = 24;
        di_im[4] = 6;
        di_re[5] = 6;
        di_im[5] = 42;
        di_re[6] = 29;
        di_im[6] = 13;
        di_re[7] = 42;
        di_im[7] = 3;
        di_re[8] = 22;
        di_im[8] = 35;
        di_re[9] = 16;
        di_im[9] = 19;
        di_re[10] = 25;
        di_im[10] = 43;
        di_re[11] = 37;
        di_im[11] = 3;
        di_re[12] = 13;
        di_im[12] = 18;
        di_re[13] = 42;
        di_im[13] = 20;
        di_re[14] = 12;
        di_im[14] = 29;
        di_re[15] = 23;
        di_im[15] = 43;

        @(posedge clk);
        di_en = 1;
        di_re[0] = 45;
        di_im[0] = 39;
        di_re[1] = 34;
        di_im[1] = 36;
        di_re[2] = 43;
        di_im[2] = 3;
        di_re[3] = 16;
        di_im[3] = 0;
        di_re[4] = 40;
        di_im[4] = 24;
        di_re[5] = 18;
        di_im[5] = 11;
        di_re[6] = 26;
        di_im[6] = 14;
        di_re[7] = 3;
        di_im[7] = 4;
        di_re[8] = 3;
        di_im[8] = 20;
        di_re[9] = 6;
        di_im[9] = 21;
        di_re[10] = 43;
        di_im[10] = 17;
        di_re[11] = 6;
        di_im[11] = 27;
        di_re[12] = 42;
        di_im[12] = 17;
        di_re[13] = 2;
        di_im[13] = 7;
        di_re[14] = 4;
        di_im[14] = 36;
        di_re[15] = 22;
        di_im[15] = 32;

        @(posedge clk);
        di_en = 1;
        di_re[0] = 34;
        di_im[0] = 27;
        di_re[1] = 30;
        di_im[1] = 42;
        di_re[2] = 32;
        di_im[2] = 42;
        di_re[3] = 22;
        di_im[3] = 7;
        di_re[4] = 3;
        di_im[4] = 34;
        di_re[5] = 15;
        di_im[5] = 32;
        di_re[6] = 31;
        di_im[6] = 25;
        di_re[7] = 34;
        di_im[7] = 24;
        di_re[8] = 23;
        di_im[8] = 24;
        di_re[9] = 45;
        di_im[9] = 19;
        di_re[10] = 6;
        di_im[10] = 12;
        di_re[11] = 33;
        di_im[11] = 40;
        di_re[12] = 47;
        di_im[12] = 10;
        di_re[13] = 36;
        di_im[13] = 28;
        di_re[14] = 19;
        di_im[14] = 24;
        di_re[15] = 24;
        di_im[15] = 31;

        @(posedge clk);
        di_en = 1;
        di_re[0] = 36;
        di_im[0] = 14;
        di_re[1] = 4;
        di_im[1] = 40;
        di_re[2] = 19;
        di_im[2] = 37;
        di_re[3] = 9;
        di_im[3] = 5;
        di_re[4] = 43;
        di_im[4] = 42;
        di_re[5] = 48;
        di_im[5] = 41;
        di_re[6] = 2;
        di_im[6] = 26;
        di_re[7] = 48;
        di_im[7] = 25;
        di_re[8] = 42;
        di_im[8] = 3;
        di_re[9] = 47;
        di_im[9] = 44;
        di_re[10] = 27;
        di_im[10] = 21;
        di_re[11] = 16;
        di_im[11] = 35;
        di_re[12] = 1;
        di_im[12] = 18;
        di_re[13] = 44;
        di_im[13] = 26;
        di_re[14] = 23;
        di_im[14] = 24;
        di_re[15] = 15;
        di_im[15] = 46;

        @(posedge clk);
        di_en = 1;
        di_re[0] = 47;
        di_im[0] = 25;
        di_re[1] = 48;
        di_im[1] = 22;
        di_re[2] = 20;
        di_im[2] = 10;
        di_re[3] = 9;
        di_im[3] = 40;
        di_re[4] = 35;
        di_im[4] = 25;
        di_re[5] = 40;
        di_im[5] = 25;
        di_re[6] = 26;
        di_im[6] = 10;
        di_re[7] = 28;
        di_im[7] = 7;
        di_re[8] = 3;
        di_im[8] = 33;
        di_re[9] = 29;
        di_im[9] = 11;
        di_re[10] = 20;
        di_im[10] = 30;
        di_re[11] = 27;
        di_im[11] = 6;
        di_re[12] = 8;
        di_im[12] = 0;
        di_re[13] = 20;
        di_im[13] = 23;
        di_re[14] = 8;
        di_im[14] = 32;
        di_re[15] = 1;
        di_im[15] = 6;

        @(posedge clk);
        di_en = 1;
        di_re[0] = 46;
        di_im[0] = 47;
        di_re[1] = 1;
        di_im[1] = 24;
        di_re[2] = 41;
        di_im[2] = 12;
        di_re[3] = 40;
        di_im[3] = 39;
        di_re[4] = 30;
        di_im[4] = 0;
        di_re[5] = 18;
        di_im[5] = 43;
        di_re[6] = 33;
        di_im[6] = 18;
        di_re[7] = 30;
        di_im[7] = 12;
        di_re[8] = 27;
        di_im[8] = 47;
        di_re[9] = 41;
        di_im[9] = 14;
        di_re[10] = 33;
        di_im[10] = 17;
        di_re[11] = 47;
        di_im[11] = 4;
        di_re[12] = 12;
        di_im[12] = 39;
        di_re[13] = 4;
        di_im[13] = 26;
        di_re[14] = 38;
        di_im[14] = 35;
        di_re[15] = 7;
        di_im[15] = 21;

        @(posedge clk);
        di_en = 1;
        di_re[0] = 17;
        di_im[0] = 23;
        di_re[1] = 28;
        di_im[1] = 7;
        di_re[2] = 43;
        di_im[2] = 31;
        di_re[3] = 8;
        di_im[3] = 27;
        di_re[4] = 45;
        di_im[4] = 38;
        di_re[5] = 33;
        di_im[5] = 22;
        di_re[6] = 12;
        di_im[6] = 27;
        di_re[7] = 12;
        di_im[7] = 15;
        di_re[8] = 44;
        di_im[8] = 42;
        di_re[9] = 38;
        di_im[9] = 44;
        di_re[10] = 9;
        di_im[10] = 25;
        di_re[11] = 30;
        di_im[11] = 44;
        di_re[12] = 32;
        di_im[12] = 19;
        di_re[13] = 36;
        di_im[13] = 39;
        di_re[14] = 29;
        di_im[14] = 4;
        di_re[15] = 44;
        di_im[15] = 3;

        @(posedge clk);
        di_en = 1;
        di_re[0] = 25;
        di_im[0] = 6;
        di_re[1] = 18;
        di_im[1] = 39;
        di_re[2] = 12;
        di_im[2] = 42;
        di_re[3] = 34;
        di_im[3] = 18;
        di_re[4] = 12;
        di_im[4] = 12;
        di_re[5] = 37;
        di_im[5] = 2;
        di_re[6] = 33;
        di_im[6] = 30;
        di_re[7] = 36;
        di_im[7] = 47;
        di_re[8] = 18;
        di_im[8] = 12;
        di_re[9] = 42;
        di_im[9] = 39;
        di_re[10] = 22;
        di_im[10] = 4;
        di_re[11] = 27;
        di_im[11] = 9;
        di_re[12] = 26;
        di_im[12] = 17;
        di_re[13] = 15;
        di_im[13] = 35;
        di_re[14] = 25;
        di_im[14] = 38;
        di_re[15] = 10;
        di_im[15] = 33;

        @(posedge clk);
        di_en = 1;
        di_re[0] = 3;
        di_im[0] = 38;
        di_re[1] = 33;
        di_im[1] = 45;
        di_re[2] = 4;
        di_im[2] = 44;
        di_re[3] = 24;
        di_im[3] = 30;
        di_re[4] = 15;
        di_im[4] = 4;
        di_re[5] = 41;
        di_im[5] = 7;
        di_re[6] = 18;
        di_im[6] = 30;
        di_re[7] = 48;
        di_im[7] = 25;
        di_re[8] = 48;
        di_im[8] = 11;
        di_re[9] = 19;
        di_im[9] = 33;
        di_re[10] = 3;
        di_im[10] = 36;
        di_re[11] = 20;
        di_im[11] = 39;
        di_re[12] = 18;
        di_im[12] = 15;
        di_re[13] = 47;
        di_im[13] = 34;
        di_re[14] = 20;
        di_im[14] = 5;
        di_re[15] = 35;
        di_im[15] = 31;

        @(posedge clk);
        di_en = 1;
        di_re[0] = 4;
        di_im[0] = 6;
        di_re[1] = 47;
        di_im[1] = 24;
        di_re[2] = 1;
        di_im[2] = 3;
        di_re[3] = 7;
        di_im[3] = 43;
        di_re[4] = 22;
        di_im[4] = 27;
        di_re[5] = 24;
        di_im[5] = 3;
        di_re[6] = 43;
        di_im[6] = 14;
        di_re[7] = 13;
        di_im[7] = 29;
        di_re[8] = 23;
        di_im[8] = 18;
        di_re[9] = 31;
        di_im[9] = 45;
        di_re[10] = 30;
        di_im[10] = 14;
        di_re[11] = 10;
        di_im[11] = 21;
        di_re[12] = 1;
        di_im[12] = 42;
        di_re[13] = 29;
        di_im[13] = 10;
        di_re[14] = 25;
        di_im[14] = 3;
        di_re[15] = 41;
        di_im[15] = 21;

        @(posedge clk);
        di_en = 1;
        di_re[0] = 26;
        di_im[0] = 27;
        di_re[1] = 33;
        di_im[1] = 18;
        di_re[2] = 4;
        di_im[2] = 22;
        di_re[3] = 2;
        di_im[3] = 35;
        di_re[4] = 2;
        di_im[4] = 46;
        di_re[5] = 36;
        di_im[5] = 45;
        di_re[6] = 25;
        di_im[6] = 12;
        di_re[7] = 12;
        di_im[7] = 36;
        di_re[8] = 48;
        di_im[8] = 17;
        di_re[9] = 36;
        di_im[9] = 5;
        di_re[10] = 29;
        di_im[10] = 21;
        di_re[11] = 35;
        di_im[11] = 13;
        di_re[12] = 5;
        di_im[12] = 22;
        di_re[13] = 31;
        di_im[13] = 6;
        di_re[14] = 22;
        di_im[14] = 31;
        di_re[15] = 40;
        di_im[15] = 15;

	@(posedge clk);
        di_en = 0;
        #3000;  // 시뮬레이션 진행 시간 확보

        $display("[TB] Simulation finished");
        $finish;
    end

    // ✅ do 출력 결과를 시뮬레이션 동안 기록

    initial begin
        fp = $fopen("do_output.txt", "w");
    end

    always @(posedge clk) begin
        for (int i = 0; i < 16; i++) begin
            $fwrite(fp, "bfly02=%0d+j%0d\n", do_re[i], do_im[i]);
        end
    end

    final begin
        $fclose(fp);
    end
endmodule

