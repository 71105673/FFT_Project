`timescale 1ns / 1ps

module tb_fft_top;

    parameter WIDTH = 9;
    parameter WIDTH_DO = 13;

    logic clk, rstn;
    logic fft_mode;
    logic di_en;
    logic signed [WIDTH-1:0] di_re[0:15];
    logic signed [WIDTH-1:0] di_im[0:15];

    logic signed [WIDTH_DO-1:0] do_re[0:15];
    logic signed [WIDTH_DO-1:0] do_im[0:15];

    integer fp;

    // // DUT
    // sdf1 #(
    //     .N(512),
    //     .M(512),
    //     .WIDTH(WIDTH),
    //     .WIDTH_DO(WIDTH_DO)
    // ) dut (
    //     .clk(clk),
    //     .rstn(rstn),
    //     .fft_mode(fft_mode),
    //     .di_en(di_en),
    //     .di_re(di_re),
    //     .di_im(di_im),

    //     .do_index(do_index),
    //     .do_en(do_en),
    //     .do_re(do_re),
    //     .do_im(do_im)
    // );

    fft_top #(
        .WIDTH(9)
    ) dut (
        .clk(clk),
        .rstn(rstn),
        .fft_mode(fft_mode),

        .din_i(di_re),
        .din_q(di_im),
        .din_valid(di_en),

        .do_re(do_re),
        .do_im(do_im),
        .do_en(do_en)
    );

    // Clock
    initial clk = 0;
    always #5 clk = ~clk;

    // Stimulus
    initial begin
        rstn = 0;
        di_en = 0;
        fft_mode = 1;
        #20;
        rstn = 1;
        #10;
        @(posedge clk);
        di_en = 1;
        di_re[0] = 63;
        di_im[0] = 0;
        di_re[1] = 64;
        di_im[1] = 0;
        di_re[2] = 64;
        di_im[2] = 0;
        di_re[3] = 64;
        di_im[3] = 0;
        di_re[4] = 64;
        di_im[4] = 0;
        di_re[5] = 64;
        di_im[5] = 0;
        di_re[6] = 64;
        di_im[6] = 0;
        di_re[7] = 64;
        di_im[7] = 0;
        di_re[8] = 64;
        di_im[8] = 0;
        di_re[9] = 64;
        di_im[9] = 0;
        di_re[10] = 64;
        di_im[10] = 0;
        di_re[11] = 63;
        di_im[11] = 0;
        di_re[12] = 63;
        di_im[12] = 0;
        di_re[13] = 63;
        di_im[13] = 0;
        di_re[14] = 63;
        di_im[14] = 0;
        di_re[15] = 63;
        di_im[15] = 0;
        @(posedge clk);
        di_en = 1;
        di_re[0] = 63;
        di_im[0] = 0;
        di_re[1] = 63;
        di_im[1] = 0;
        di_re[2] = 62;
        di_im[2] = 0;
        di_re[3] = 62;
        di_im[3] = 0;
        di_re[4] = 62;
        di_im[4] = 0;
        di_re[5] = 62;
        di_im[5] = 0;
        di_re[6] = 62;
        di_im[6] = 0;
        di_re[7] = 61;
        di_im[7] = 0;
        di_re[8] = 61;
        di_im[8] = 0;
        di_re[9] = 61;
        di_im[9] = 0;
        di_re[10] = 61;
        di_im[10] = 0;
        di_re[11] = 61;
        di_im[11] = 0;
        di_re[12] = 60;
        di_im[12] = 0;
        di_re[13] = 60;
        di_im[13] = 0;
        di_re[14] = 60;
        di_im[14] = 0;
        di_re[15] = 59;
        di_im[15] = 0;
        @(posedge clk);
        di_en = 1;
        di_re[0] = 59;
        di_im[0] = 0;
        di_re[1] = 59;
        di_im[1] = 0;
        di_re[2] = 59;
        di_im[2] = 0;
        di_re[3] = 58;
        di_im[3] = 0;
        di_re[4] = 58;
        di_im[4] = 0;
        di_re[5] = 58;
        di_im[5] = 0;
        di_re[6] = 57;
        di_im[6] = 0;
        di_re[7] = 57;
        di_im[7] = 0;
        di_re[8] = 56;
        di_im[8] = 0;
        di_re[9] = 56;
        di_im[9] = 0;
        di_re[10] = 56;
        di_im[10] = 0;
        di_re[11] = 55;
        di_im[11] = 0;
        di_re[12] = 55;
        di_im[12] = 0;
        di_re[13] = 54;
        di_im[13] = 0;
        di_re[14] = 54;
        di_im[14] = 0;
        di_re[15] = 54;
        di_im[15] = 0;
        @(posedge clk);
        di_en = 1;
        di_re[0] = 53;
        di_im[0] = 0;
        di_re[1] = 53;
        di_im[1] = 0;
        di_re[2] = 52;
        di_im[2] = 0;
        di_re[3] = 52;
        di_im[3] = 0;
        di_re[4] = 51;
        di_im[4] = 0;
        di_re[5] = 51;
        di_im[5] = 0;
        di_re[6] = 50;
        di_im[6] = 0;
        di_re[7] = 50;
        di_im[7] = 0;
        di_re[8] = 49;
        di_im[8] = 0;
        di_re[9] = 49;
        di_im[9] = 0;
        di_re[10] = 48;
        di_im[10] = 0;
        di_re[11] = 48;
        di_im[11] = 0;
        di_re[12] = 47;
        di_im[12] = 0;
        di_re[13] = 47;
        di_im[13] = 0;
        di_re[14] = 46;
        di_im[14] = 0;
        di_re[15] = 46;
        di_im[15] = 0;
        @(posedge clk);
        di_en = 1;
        di_re[0] = 45;
        di_im[0] = 0;
        di_re[1] = 45;
        di_im[1] = 0;
        di_re[2] = 44;
        di_im[2] = 0;
        di_re[3] = 44;
        di_im[3] = 0;
        di_re[4] = 43;
        di_im[4] = 0;
        di_re[5] = 42;
        di_im[5] = 0;
        di_re[6] = 42;
        di_im[6] = 0;
        di_re[7] = 41;
        di_im[7] = 0;
        di_re[8] = 41;
        di_im[8] = 0;
        di_re[9] = 40;
        di_im[9] = 0;
        di_re[10] = 39;
        di_im[10] = 0;
        di_re[11] = 39;
        di_im[11] = 0;
        di_re[12] = 38;
        di_im[12] = 0;
        di_re[13] = 37;
        di_im[13] = 0;
        di_re[14] = 37;
        di_im[14] = 0;
        di_re[15] = 36;
        di_im[15] = 0;
        @(posedge clk);
        di_en = 1;
        di_re[0] = 36;
        di_im[0] = 0;
        di_re[1] = 35;
        di_im[1] = 0;
        di_re[2] = 34;
        di_im[2] = 0;
        di_re[3] = 34;
        di_im[3] = 0;
        di_re[4] = 33;
        di_im[4] = 0;
        di_re[5] = 32;
        di_im[5] = 0;
        di_re[6] = 32;
        di_im[6] = 0;
        di_re[7] = 31;
        di_im[7] = 0;
        di_re[8] = 30;
        di_im[8] = 0;
        di_re[9] = 29;
        di_im[9] = 0;
        di_re[10] = 29;
        di_im[10] = 0;
        di_re[11] = 28;
        di_im[11] = 0;
        di_re[12] = 27;
        di_im[12] = 0;
        di_re[13] = 27;
        di_im[13] = 0;
        di_re[14] = 26;
        di_im[14] = 0;
        di_re[15] = 25;
        di_im[15] = 0;
        @(posedge clk);
        di_en = 1;
        di_re[0] = 24;
        di_im[0] = 0;
        di_re[1] = 24;
        di_im[1] = 0;
        di_re[2] = 23;
        di_im[2] = 0;
        di_re[3] = 22;
        di_im[3] = 0;
        di_re[4] = 22;
        di_im[4] = 0;
        di_re[5] = 21;
        di_im[5] = 0;
        di_re[6] = 20;
        di_im[6] = 0;
        di_re[7] = 19;
        di_im[7] = 0;
        di_re[8] = 19;
        di_im[8] = 0;
        di_re[9] = 18;
        di_im[9] = 0;
        di_re[10] = 17;
        di_im[10] = 0;
        di_re[11] = 16;
        di_im[11] = 0;
        di_re[12] = 16;
        di_im[12] = 0;
        di_re[13] = 15;
        di_im[13] = 0;
        di_re[14] = 14;
        di_im[14] = 0;
        di_re[15] = 13;
        di_im[15] = 0;
        @(posedge clk);
        di_en = 1;
        di_re[0] = 12;
        di_im[0] = 0;
        di_re[1] = 12;
        di_im[1] = 0;
        di_re[2] = 11;
        di_im[2] = 0;
        di_re[3] = 10;
        di_im[3] = 0;
        di_re[4] = 9;
        di_im[4] = 0;
        di_re[5] = 9;
        di_im[5] = 0;
        di_re[6] = 8;
        di_im[6] = 0;
        di_re[7] = 7;
        di_im[7] = 0;
        di_re[8] = 6;
        di_im[8] = 0;
        di_re[9] = 5;
        di_im[9] = 0;
        di_re[10] = 5;
        di_im[10] = 0;
        di_re[11] = 4;
        di_im[11] = 0;
        di_re[12] = 3;
        di_im[12] = 0;
        di_re[13] = 2;
        di_im[13] = 0;
        di_re[14] = 2;
        di_im[14] = 0;
        di_re[15] = 1;
        di_im[15] = 0;
        @(posedge clk);
        di_en = 1;
        di_re[0] = 0;
        di_im[0] = 0;
        di_re[1] = -1;
        di_im[1] = 0;
        di_re[2] = -2;
        di_im[2] = 0;
        di_re[3] = -2;
        di_im[3] = 0;
        di_re[4] = -3;
        di_im[4] = 0;
        di_re[5] = -4;
        di_im[5] = 0;
        di_re[6] = -5;
        di_im[6] = 0;
        di_re[7] = -5;
        di_im[7] = 0;
        di_re[8] = -6;
        di_im[8] = 0;
        di_re[9] = -7;
        di_im[9] = 0;
        di_re[10] = -8;
        di_im[10] = 0;
        di_re[11] = -9;
        di_im[11] = 0;
        di_re[12] = -9;
        di_im[12] = 0;
        di_re[13] = -10;
        di_im[13] = 0;
        di_re[14] = -11;
        di_im[14] = 0;
        di_re[15] = -12;
        di_im[15] = 0;
        @(posedge clk);
        di_en = 1;
        di_re[0] = -12;
        di_im[0] = 0;
        di_re[1] = -13;
        di_im[1] = 0;
        di_re[2] = -14;
        di_im[2] = 0;
        di_re[3] = -15;
        di_im[3] = 0;
        di_re[4] = -16;
        di_im[4] = 0;
        di_re[5] = -16;
        di_im[5] = 0;
        di_re[6] = -17;
        di_im[6] = 0;
        di_re[7] = -18;
        di_im[7] = 0;
        di_re[8] = -19;
        di_im[8] = 0;
        di_re[9] = -19;
        di_im[9] = 0;
        di_re[10] = -20;
        di_im[10] = 0;
        di_re[11] = -21;
        di_im[11] = 0;
        di_re[12] = -22;
        di_im[12] = 0;
        di_re[13] = -22;
        di_im[13] = 0;
        di_re[14] = -23;
        di_im[14] = 0;
        di_re[15] = -24;
        di_im[15] = 0;
        @(posedge clk);
        di_en = 1;
        di_re[0] = -24;
        di_im[0] = 0;
        di_re[1] = -25;
        di_im[1] = 0;
        di_re[2] = -26;
        di_im[2] = 0;
        di_re[3] = -27;
        di_im[3] = 0;
        di_re[4] = -27;
        di_im[4] = 0;
        di_re[5] = -28;
        di_im[5] = 0;
        di_re[6] = -29;
        di_im[6] = 0;
        di_re[7] = -29;
        di_im[7] = 0;
        di_re[8] = -30;
        di_im[8] = 0;
        di_re[9] = -31;
        di_im[9] = 0;
        di_re[10] = -32;
        di_im[10] = 0;
        di_re[11] = -32;
        di_im[11] = 0;
        di_re[12] = -33;
        di_im[12] = 0;
        di_re[13] = -34;
        di_im[13] = 0;
        di_re[14] = -34;
        di_im[14] = 0;
        di_re[15] = -35;
        di_im[15] = 0;
        @(posedge clk);
        di_en = 1;
        di_re[0] = -36;
        di_im[0] = 0;
        di_re[1] = -36;
        di_im[1] = 0;
        di_re[2] = -37;
        di_im[2] = 0;
        di_re[3] = -37;
        di_im[3] = 0;
        di_re[4] = -38;
        di_im[4] = 0;
        di_re[5] = -39;
        di_im[5] = 0;
        di_re[6] = -39;
        di_im[6] = 0;
        di_re[7] = -40;
        di_im[7] = 0;
        di_re[8] = -41;
        di_im[8] = 0;
        di_re[9] = -41;
        di_im[9] = 0;
        di_re[10] = -42;
        di_im[10] = 0;
        di_re[11] = -42;
        di_im[11] = 0;
        di_re[12] = -43;
        di_im[12] = 0;
        di_re[13] = -44;
        di_im[13] = 0;
        di_re[14] = -44;
        di_im[14] = 0;
        di_re[15] = -45;
        di_im[15] = 0;
        @(posedge clk);
        di_en = 1;
        di_re[0] = -45;
        di_im[0] = 0;
        di_re[1] = -46;
        di_im[1] = 0;
        di_re[2] = -46;
        di_im[2] = 0;
        di_re[3] = -47;
        di_im[3] = 0;
        di_re[4] = -47;
        di_im[4] = 0;
        di_re[5] = -48;
        di_im[5] = 0;
        di_re[6] = -48;
        di_im[6] = 0;
        di_re[7] = -49;
        di_im[7] = 0;
        di_re[8] = -49;
        di_im[8] = 0;
        di_re[9] = -50;
        di_im[9] = 0;
        di_re[10] = -50;
        di_im[10] = 0;
        di_re[11] = -51;
        di_im[11] = 0;
        di_re[12] = -51;
        di_im[12] = 0;
        di_re[13] = -52;
        di_im[13] = 0;
        di_re[14] = -52;
        di_im[14] = 0;
        di_re[15] = -53;
        di_im[15] = 0;
        @(posedge clk);
        di_en = 1;
        di_re[0] = -53;
        di_im[0] = 0;
        di_re[1] = -54;
        di_im[1] = 0;
        di_re[2] = -54;
        di_im[2] = 0;
        di_re[3] = -54;
        di_im[3] = 0;
        di_re[4] = -55;
        di_im[4] = 0;
        di_re[5] = -55;
        di_im[5] = 0;
        di_re[6] = -56;
        di_im[6] = 0;
        di_re[7] = -56;
        di_im[7] = 0;
        di_re[8] = -56;
        di_im[8] = 0;
        di_re[9] = -57;
        di_im[9] = 0;
        di_re[10] = -57;
        di_im[10] = 0;
        di_re[11] = -58;
        di_im[11] = 0;
        di_re[12] = -58;
        di_im[12] = 0;
        di_re[13] = -58;
        di_im[13] = 0;
        di_re[14] = -59;
        di_im[14] = 0;
        di_re[15] = -59;
        di_im[15] = 0;
        @(posedge clk);
        di_en = 1;
        di_re[0] = -59;
        di_im[0] = 0;
        di_re[1] = -59;
        di_im[1] = 0;
        di_re[2] = -60;
        di_im[2] = 0;
        di_re[3] = -60;
        di_im[3] = 0;
        di_re[4] = -60;
        di_im[4] = 0;
        di_re[5] = -61;
        di_im[5] = 0;
        di_re[6] = -61;
        di_im[6] = 0;
        di_re[7] = -61;
        di_im[7] = 0;
        di_re[8] = -61;
        di_im[8] = 0;
        di_re[9] = -61;
        di_im[9] = 0;
        di_re[10] = -62;
        di_im[10] = 0;
        di_re[11] = -62;
        di_im[11] = 0;
        di_re[12] = -62;
        di_im[12] = 0;
        di_re[13] = -62;
        di_im[13] = 0;
        di_re[14] = -62;
        di_im[14] = 0;
        di_re[15] = -63;
        di_im[15] = 0;
        @(posedge clk);
        di_en = 1;
        di_re[0] = -63;
        di_im[0] = 0;
        di_re[1] = -63;
        di_im[1] = 0;
        di_re[2] = -63;
        di_im[2] = 0;
        di_re[3] = -63;
        di_im[3] = 0;
        di_re[4] = -63;
        di_im[4] = 0;
        di_re[5] = -63;
        di_im[5] = 0;
        di_re[6] = -64;
        di_im[6] = 0;
        di_re[7] = -64;
        di_im[7] = 0;
        di_re[8] = -64;
        di_im[8] = 0;
        di_re[9] = -64;
        di_im[9] = 0;
        di_re[10] = -64;
        di_im[10] = 0;
        di_re[11] = -64;
        di_im[11] = 0;
        di_re[12] = -64;
        di_im[12] = 0;
        di_re[13] = -64;
        di_im[13] = 0;
        di_re[14] = -64;
        di_im[14] = 0;
        di_re[15] = -64;
        di_im[15] = 0;
        @(posedge clk);
        di_en = 1;
        di_re[0] = -64;
        di_im[0] = 0;
        di_re[1] = -64;
        di_im[1] = 0;
        di_re[2] = -64;
        di_im[2] = 0;
        di_re[3] = -64;
        di_im[3] = 0;
        di_re[4] = -64;
        di_im[4] = 0;
        di_re[5] = -64;
        di_im[5] = 0;
        di_re[6] = -64;
        di_im[6] = 0;
        di_re[7] = -64;
        di_im[7] = 0;
        di_re[8] = -64;
        di_im[8] = 0;
        di_re[9] = -64;
        di_im[9] = 0;
        di_re[10] = -64;
        di_im[10] = 0;
        di_re[11] = -63;
        di_im[11] = 0;
        di_re[12] = -63;
        di_im[12] = 0;
        di_re[13] = -63;
        di_im[13] = 0;
        di_re[14] = -63;
        di_im[14] = 0;
        di_re[15] = -63;
        di_im[15] = 0;
        @(posedge clk);
        di_en = 1;
        di_re[0] = -63;
        di_im[0] = 0;
        di_re[1] = -63;
        di_im[1] = 0;
        di_re[2] = -62;
        di_im[2] = 0;
        di_re[3] = -62;
        di_im[3] = 0;
        di_re[4] = -62;
        di_im[4] = 0;
        di_re[5] = -62;
        di_im[5] = 0;
        di_re[6] = -62;
        di_im[6] = 0;
        di_re[7] = -61;
        di_im[7] = 0;
        di_re[8] = -61;
        di_im[8] = 0;
        di_re[9] = -61;
        di_im[9] = 0;
        di_re[10] = -61;
        di_im[10] = 0;
        di_re[11] = -61;
        di_im[11] = 0;
        di_re[12] = -60;
        di_im[12] = 0;
        di_re[13] = -60;
        di_im[13] = 0;
        di_re[14] = -60;
        di_im[14] = 0;
        di_re[15] = -59;
        di_im[15] = 0;
        @(posedge clk);
        di_en = 1;
        di_re[0] = -59;
        di_im[0] = 0;
        di_re[1] = -59;
        di_im[1] = 0;
        di_re[2] = -59;
        di_im[2] = 0;
        di_re[3] = -58;
        di_im[3] = 0;
        di_re[4] = -58;
        di_im[4] = 0;
        di_re[5] = -58;
        di_im[5] = 0;
        di_re[6] = -57;
        di_im[6] = 0;
        di_re[7] = -57;
        di_im[7] = 0;
        di_re[8] = -56;
        di_im[8] = 0;
        di_re[9] = -56;
        di_im[9] = 0;
        di_re[10] = -56;
        di_im[10] = 0;
        di_re[11] = -55;
        di_im[11] = 0;
        di_re[12] = -55;
        di_im[12] = 0;
        di_re[13] = -54;
        di_im[13] = 0;
        di_re[14] = -54;
        di_im[14] = 0;
        di_re[15] = -54;
        di_im[15] = 0;
        @(posedge clk);
        di_en = 1;
        di_re[0] = -53;
        di_im[0] = 0;
        di_re[1] = -53;
        di_im[1] = 0;
        di_re[2] = -52;
        di_im[2] = 0;
        di_re[3] = -52;
        di_im[3] = 0;
        di_re[4] = -51;
        di_im[4] = 0;
        di_re[5] = -51;
        di_im[5] = 0;
        di_re[6] = -50;
        di_im[6] = 0;
        di_re[7] = -50;
        di_im[7] = 0;
        di_re[8] = -49;
        di_im[8] = 0;
        di_re[9] = -49;
        di_im[9] = 0;
        di_re[10] = -48;
        di_im[10] = 0;
        di_re[11] = -48;
        di_im[11] = 0;
        di_re[12] = -47;
        di_im[12] = 0;
        di_re[13] = -47;
        di_im[13] = 0;
        di_re[14] = -46;
        di_im[14] = 0;
        di_re[15] = -46;
        di_im[15] = 0;
        @(posedge clk);
        di_en = 1;
        di_re[0] = -45;
        di_im[0] = 0;
        di_re[1] = -45;
        di_im[1] = 0;
        di_re[2] = -44;
        di_im[2] = 0;
        di_re[3] = -44;
        di_im[3] = 0;
        di_re[4] = -43;
        di_im[4] = 0;
        di_re[5] = -42;
        di_im[5] = 0;
        di_re[6] = -42;
        di_im[6] = 0;
        di_re[7] = -41;
        di_im[7] = 0;
        di_re[8] = -41;
        di_im[8] = 0;
        di_re[9] = -40;
        di_im[9] = 0;
        di_re[10] = -39;
        di_im[10] = 0;
        di_re[11] = -39;
        di_im[11] = 0;
        di_re[12] = -38;
        di_im[12] = 0;
        di_re[13] = -37;
        di_im[13] = 0;
        di_re[14] = -37;
        di_im[14] = 0;
        di_re[15] = -36;
        di_im[15] = 0;
        @(posedge clk);
        di_en = 1;
        di_re[0] = -36;
        di_im[0] = 0;
        di_re[1] = -35;
        di_im[1] = 0;
        di_re[2] = -34;
        di_im[2] = 0;
        di_re[3] = -34;
        di_im[3] = 0;
        di_re[4] = -33;
        di_im[4] = 0;
        di_re[5] = -32;
        di_im[5] = 0;
        di_re[6] = -32;
        di_im[6] = 0;
        di_re[7] = -31;
        di_im[7] = 0;
        di_re[8] = -30;
        di_im[8] = 0;
        di_re[9] = -29;
        di_im[9] = 0;
        di_re[10] = -29;
        di_im[10] = 0;
        di_re[11] = -28;
        di_im[11] = 0;
        di_re[12] = -27;
        di_im[12] = 0;
        di_re[13] = -27;
        di_im[13] = 0;
        di_re[14] = -26;
        di_im[14] = 0;
        di_re[15] = -25;
        di_im[15] = 0;
        @(posedge clk);
        di_en = 1;
        di_re[0] = -24;
        di_im[0] = 0;
        di_re[1] = -24;
        di_im[1] = 0;
        di_re[2] = -23;
        di_im[2] = 0;
        di_re[3] = -22;
        di_im[3] = 0;
        di_re[4] = -22;
        di_im[4] = 0;
        di_re[5] = -21;
        di_im[5] = 0;
        di_re[6] = -20;
        di_im[6] = 0;
        di_re[7] = -19;
        di_im[7] = 0;
        di_re[8] = -19;
        di_im[8] = 0;
        di_re[9] = -18;
        di_im[9] = 0;
        di_re[10] = -17;
        di_im[10] = 0;
        di_re[11] = -16;
        di_im[11] = 0;
        di_re[12] = -16;
        di_im[12] = 0;
        di_re[13] = -15;
        di_im[13] = 0;
        di_re[14] = -14;
        di_im[14] = 0;
        di_re[15] = -13;
        di_im[15] = 0;
        @(posedge clk);
        di_en = 1;
        di_re[0] = -12;
        di_im[0] = 0;
        di_re[1] = -12;
        di_im[1] = 0;
        di_re[2] = -11;
        di_im[2] = 0;
        di_re[3] = -10;
        di_im[3] = 0;
        di_re[4] = -9;
        di_im[4] = 0;
        di_re[5] = -9;
        di_im[5] = 0;
        di_re[6] = -8;
        di_im[6] = 0;
        di_re[7] = -7;
        di_im[7] = 0;
        di_re[8] = -6;
        di_im[8] = 0;
        di_re[9] = -5;
        di_im[9] = 0;
        di_re[10] = -5;
        di_im[10] = 0;
        di_re[11] = -4;
        di_im[11] = 0;
        di_re[12] = -3;
        di_im[12] = 0;
        di_re[13] = -2;
        di_im[13] = 0;
        di_re[14] = -2;
        di_im[14] = 0;
        di_re[15] = -1;
        di_im[15] = 0;
        @(posedge clk);
        di_en = 1;
        di_re[0] = 0;
        di_im[0] = 0;
        di_re[1] = 1;
        di_im[1] = 0;
        di_re[2] = 2;
        di_im[2] = 0;
        di_re[3] = 2;
        di_im[3] = 0;
        di_re[4] = 3;
        di_im[4] = 0;
        di_re[5] = 4;
        di_im[5] = 0;
        di_re[6] = 5;
        di_im[6] = 0;
        di_re[7] = 5;
        di_im[7] = 0;
        di_re[8] = 6;
        di_im[8] = 0;
        di_re[9] = 7;
        di_im[9] = 0;
        di_re[10] = 8;
        di_im[10] = 0;
        di_re[11] = 9;
        di_im[11] = 0;
        di_re[12] = 9;
        di_im[12] = 0;
        di_re[13] = 10;
        di_im[13] = 0;
        di_re[14] = 11;
        di_im[14] = 0;
        di_re[15] = 12;
        di_im[15] = 0;
        @(posedge clk);
        di_en = 1;
        di_re[0] = 12;
        di_im[0] = 0;
        di_re[1] = 13;
        di_im[1] = 0;
        di_re[2] = 14;
        di_im[2] = 0;
        di_re[3] = 15;
        di_im[3] = 0;
        di_re[4] = 16;
        di_im[4] = 0;
        di_re[5] = 16;
        di_im[5] = 0;
        di_re[6] = 17;
        di_im[6] = 0;
        di_re[7] = 18;
        di_im[7] = 0;
        di_re[8] = 19;
        di_im[8] = 0;
        di_re[9] = 19;
        di_im[9] = 0;
        di_re[10] = 20;
        di_im[10] = 0;
        di_re[11] = 21;
        di_im[11] = 0;
        di_re[12] = 22;
        di_im[12] = 0;
        di_re[13] = 22;
        di_im[13] = 0;
        di_re[14] = 23;
        di_im[14] = 0;
        di_re[15] = 24;
        di_im[15] = 0;
        @(posedge clk);
        di_en = 1;
        di_re[0] = 24;
        di_im[0] = 0;
        di_re[1] = 25;
        di_im[1] = 0;
        di_re[2] = 26;
        di_im[2] = 0;
        di_re[3] = 27;
        di_im[3] = 0;
        di_re[4] = 27;
        di_im[4] = 0;
        di_re[5] = 28;
        di_im[5] = 0;
        di_re[6] = 29;
        di_im[6] = 0;
        di_re[7] = 29;
        di_im[7] = 0;
        di_re[8] = 30;
        di_im[8] = 0;
        di_re[9] = 31;
        di_im[9] = 0;
        di_re[10] = 32;
        di_im[10] = 0;
        di_re[11] = 32;
        di_im[11] = 0;
        di_re[12] = 33;
        di_im[12] = 0;
        di_re[13] = 34;
        di_im[13] = 0;
        di_re[14] = 34;
        di_im[14] = 0;
        di_re[15] = 35;
        di_im[15] = 0;
        @(posedge clk);
        di_en = 1;
        di_re[0] = 36;
        di_im[0] = 0;
        di_re[1] = 36;
        di_im[1] = 0;
        di_re[2] = 37;
        di_im[2] = 0;
        di_re[3] = 37;
        di_im[3] = 0;
        di_re[4] = 38;
        di_im[4] = 0;
        di_re[5] = 39;
        di_im[5] = 0;
        di_re[6] = 39;
        di_im[6] = 0;
        di_re[7] = 40;
        di_im[7] = 0;
        di_re[8] = 41;
        di_im[8] = 0;
        di_re[9] = 41;
        di_im[9] = 0;
        di_re[10] = 42;
        di_im[10] = 0;
        di_re[11] = 42;
        di_im[11] = 0;
        di_re[12] = 43;
        di_im[12] = 0;
        di_re[13] = 44;
        di_im[13] = 0;
        di_re[14] = 44;
        di_im[14] = 0;
        di_re[15] = 45;
        di_im[15] = 0;
        @(posedge clk);
        di_en = 1;
        di_re[0] = 45;
        di_im[0] = 0;
        di_re[1] = 46;
        di_im[1] = 0;
        di_re[2] = 46;
        di_im[2] = 0;
        di_re[3] = 47;
        di_im[3] = 0;
        di_re[4] = 47;
        di_im[4] = 0;
        di_re[5] = 48;
        di_im[5] = 0;
        di_re[6] = 48;
        di_im[6] = 0;
        di_re[7] = 49;
        di_im[7] = 0;
        di_re[8] = 49;
        di_im[8] = 0;
        di_re[9] = 50;
        di_im[9] = 0;
        di_re[10] = 50;
        di_im[10] = 0;
        di_re[11] = 51;
        di_im[11] = 0;
        di_re[12] = 51;
        di_im[12] = 0;
        di_re[13] = 52;
        di_im[13] = 0;
        di_re[14] = 52;
        di_im[14] = 0;
        di_re[15] = 53;
        di_im[15] = 0;
        @(posedge clk);
        di_en = 1;
        di_re[0] = 53;
        di_im[0] = 0;
        di_re[1] = 54;
        di_im[1] = 0;
        di_re[2] = 54;
        di_im[2] = 0;
        di_re[3] = 54;
        di_im[3] = 0;
        di_re[4] = 55;
        di_im[4] = 0;
        di_re[5] = 55;
        di_im[5] = 0;
        di_re[6] = 56;
        di_im[6] = 0;
        di_re[7] = 56;
        di_im[7] = 0;
        di_re[8] = 56;
        di_im[8] = 0;
        di_re[9] = 57;
        di_im[9] = 0;
        di_re[10] = 57;
        di_im[10] = 0;
        di_re[11] = 58;
        di_im[11] = 0;
        di_re[12] = 58;
        di_im[12] = 0;
        di_re[13] = 58;
        di_im[13] = 0;
        di_re[14] = 59;
        di_im[14] = 0;
        di_re[15] = 59;
        di_im[15] = 0;
        @(posedge clk);
        di_en = 1;
        di_re[0] = 59;
        di_im[0] = 0;
        di_re[1] = 59;
        di_im[1] = 0;
        di_re[2] = 60;
        di_im[2] = 0;
        di_re[3] = 60;
        di_im[3] = 0;
        di_re[4] = 60;
        di_im[4] = 0;
        di_re[5] = 61;
        di_im[5] = 0;
        di_re[6] = 61;
        di_im[6] = 0;
        di_re[7] = 61;
        di_im[7] = 0;
        di_re[8] = 61;
        di_im[8] = 0;
        di_re[9] = 61;
        di_im[9] = 0;
        di_re[10] = 62;
        di_im[10] = 0;
        di_re[11] = 62;
        di_im[11] = 0;
        di_re[12] = 62;
        di_im[12] = 0;
        di_re[13] = 62;
        di_im[13] = 0;
        di_re[14] = 62;
        di_im[14] = 0;
        di_re[15] = 63;
        di_im[15] = 0;
        @(posedge clk);
        di_en = 1;
        di_re[0] = 63;
        di_im[0] = 0;
        di_re[1] = 63;
        di_im[1] = 0;
        di_re[2] = 63;
        di_im[2] = 0;
        di_re[3] = 63;
        di_im[3] = 0;
        di_re[4] = 63;
        di_im[4] = 0;
        di_re[5] = 63;
        di_im[5] = 0;
        di_re[6] = 64;
        di_im[6] = 0;
        di_re[7] = 64;
        di_im[7] = 0;
        di_re[8] = 64;
        di_im[8] = 0;
        di_re[9] = 64;
        di_im[9] = 0;
        di_re[10] = 64;
        di_im[10] = 0;
        di_re[11] = 64;
        di_im[11] = 0;
        di_re[12] = 64;
        di_im[12] = 0;
        di_re[13] = 64;
        di_im[13] = 0;
        di_re[14] = 64;
        di_im[14] = 0;
        di_re[15] = 64;
        di_im[15] = 0;
        @(posedge clk);
        di_en = 0;
        #3000;  // 시뮬레이션 진행 시간 확보

        $display("[TB] Simulation finished");
        $finish;
    end

    // ✅ do 출력 결과를 시뮬레이션 동안 기록

    initial begin
        fp = $fopen("do_output.txt", "w");
    end

    always @(posedge clk) begin
        for (int i = 0; i < 16; i++) begin
            $fwrite(fp, "bfly02=%0d+j%0d\n", do_re[i], do_im[i]);
        end
    end

    final begin
        $fclose(fp);
    end
endmodule

