`timescale 1ns / 1ps

module twiddle_512 #(
    parameter WIDTH = 9,
    parameter TW_TABLE_DEPTH = 512,
    parameter TW_FF = 1,
    parameter NUM_PARALLEL_PATHS = 16 // 이 파라미터를 추가
)(
    input clk,
    // addr를 배열로 변경: [0:NUM_PARALLEL_PATHS-1] 형태로 선언
    input [$clog2(TW_TABLE_DEPTH)-1:0] addr, 
    
    output signed [WIDTH-1:0] tw_re,
    output signed [WIDTH-1:0] tw_im
);

    wire[8:0]  twf_m0_real_val[0:TW_TABLE_DEPTH-1];   //  Twiddle Table (Real)
    wire[8:0]  twf_m0_imag_val[0:TW_TABLE_DEPTH-1];   //  Twiddle Table (Imag)
    wire[8:0]  mx_re;          //  Multiplexer output (Real)
    wire[8:0]  mx_im;          //  Multiplexer output (Imag)
    reg [8:0]  ff_re;          //  Register output (Real)
    reg [8:0]  ff_im;          //  Register output (Imag)

    assign  mx_re = twf_m0_real_val[addr];
    assign  mx_im = twf_m0_imag_val[addr];

    always @(posedge clk) begin
        ff_re <= mx_re;
        ff_im <= mx_im;
    end

    assign  tw_re = TW_FF ? ff_re : mx_re;
    assign  tw_im = TW_FF ? ff_im : mx_im;

    //----------------------------------------------------------------------
    //  Twiddle Factor Value
    //----------------------------------------------------------------------
    assign twf_m0_real_val[  0] = 9'sd128; assign twf_m0_imag_val[  0] = 9'sd0;
    assign twf_m0_real_val[  1] = 9'sd128; assign twf_m0_imag_val[  1] = 9'sd0;
    assign twf_m0_real_val[  2] = 9'sd128; assign twf_m0_imag_val[  2] = 9'sd0;
    assign twf_m0_real_val[  3] = 9'sd128; assign twf_m0_imag_val[  3] = 9'sd0;
    assign twf_m0_real_val[  4] = 9'sd128; assign twf_m0_imag_val[  4] = 9'sd0;
    assign twf_m0_real_val[  5] = 9'sd128; assign twf_m0_imag_val[  5] = 9'sd0;
    assign twf_m0_real_val[  6] = 9'sd128; assign twf_m0_imag_val[  6] = 9'sd0;
    assign twf_m0_real_val[  7] = 9'sd128; assign twf_m0_imag_val[  7] = 9'sd0;
    assign twf_m0_real_val[  8] = 9'sd128; assign twf_m0_imag_val[  8] = 9'sd0;
    assign twf_m0_real_val[  9] = 9'sd128; assign twf_m0_imag_val[  9] = 9'sd0;
    assign twf_m0_real_val[ 10] = 9'sd128; assign twf_m0_imag_val[ 10] = 9'sd0;
    assign twf_m0_real_val[ 11] = 9'sd128; assign twf_m0_imag_val[ 11] = 9'sd0;
    assign twf_m0_real_val[ 12] = 9'sd128; assign twf_m0_imag_val[ 12] = 9'sd0;
    assign twf_m0_real_val[ 13] = 9'sd128; assign twf_m0_imag_val[ 13] = 9'sd0;
    assign twf_m0_real_val[ 14] = 9'sd128; assign twf_m0_imag_val[ 14] = 9'sd0;
    assign twf_m0_real_val[ 15] = 9'sd128; assign twf_m0_imag_val[ 15] = 9'sd0;
    assign twf_m0_real_val[ 16] = 9'sd128; assign twf_m0_imag_val[ 16] = 9'sd0;
    assign twf_m0_real_val[ 17] = 9'sd128; assign twf_m0_imag_val[ 17] = 9'sd0;
    assign twf_m0_real_val[ 18] = 9'sd128; assign twf_m0_imag_val[ 18] = 9'sd0;
    assign twf_m0_real_val[ 19] = 9'sd128; assign twf_m0_imag_val[ 19] = 9'sd0;
    assign twf_m0_real_val[ 20] = 9'sd128; assign twf_m0_imag_val[ 20] = 9'sd0;
    assign twf_m0_real_val[ 21] = 9'sd128; assign twf_m0_imag_val[ 21] = 9'sd0;
    assign twf_m0_real_val[ 22] = 9'sd128; assign twf_m0_imag_val[ 22] = 9'sd0;
    assign twf_m0_real_val[ 23] = 9'sd128; assign twf_m0_imag_val[ 23] = 9'sd0;
    assign twf_m0_real_val[ 24] = 9'sd128; assign twf_m0_imag_val[ 24] = 9'sd0;
    assign twf_m0_real_val[ 25] = 9'sd128; assign twf_m0_imag_val[ 25] = 9'sd0;
    assign twf_m0_real_val[ 26] = 9'sd128; assign twf_m0_imag_val[ 26] = 9'sd0;
    assign twf_m0_real_val[ 27] = 9'sd128; assign twf_m0_imag_val[ 27] = 9'sd0;
    assign twf_m0_real_val[ 28] = 9'sd128; assign twf_m0_imag_val[ 28] = 9'sd0;
    assign twf_m0_real_val[ 29] = 9'sd128; assign twf_m0_imag_val[ 29] = 9'sd0;
    assign twf_m0_real_val[ 30] = 9'sd128; assign twf_m0_imag_val[ 30] = 9'sd0;
    assign twf_m0_real_val[ 31] = 9'sd128; assign twf_m0_imag_val[ 31] = 9'sd0;
    assign twf_m0_real_val[ 32] = 9'sd128; assign twf_m0_imag_val[ 32] = 9'sd0;
    assign twf_m0_real_val[ 33] = 9'sd128; assign twf_m0_imag_val[ 33] = 9'sd0;
    assign twf_m0_real_val[ 34] = 9'sd128; assign twf_m0_imag_val[ 34] = 9'sd0;
    assign twf_m0_real_val[ 35] = 9'sd128; assign twf_m0_imag_val[ 35] = 9'sd0;
    assign twf_m0_real_val[ 36] = 9'sd128; assign twf_m0_imag_val[ 36] = 9'sd0;
    assign twf_m0_real_val[ 37] = 9'sd128; assign twf_m0_imag_val[ 37] = 9'sd0;
    assign twf_m0_real_val[ 38] = 9'sd128; assign twf_m0_imag_val[ 38] = 9'sd0;
    assign twf_m0_real_val[ 39] = 9'sd128; assign twf_m0_imag_val[ 39] = 9'sd0;
    assign twf_m0_real_val[ 40] = 9'sd128; assign twf_m0_imag_val[ 40] = 9'sd0;
    assign twf_m0_real_val[ 41] = 9'sd128; assign twf_m0_imag_val[ 41] = 9'sd0;
    assign twf_m0_real_val[ 42] = 9'sd128; assign twf_m0_imag_val[ 42] = 9'sd0;
    assign twf_m0_real_val[ 43] = 9'sd128; assign twf_m0_imag_val[ 43] = 9'sd0;
    assign twf_m0_real_val[ 44] = 9'sd128; assign twf_m0_imag_val[ 44] = 9'sd0;
    assign twf_m0_real_val[ 45] = 9'sd128; assign twf_m0_imag_val[ 45] = 9'sd0;
    assign twf_m0_real_val[ 46] = 9'sd128; assign twf_m0_imag_val[ 46] = 9'sd0;
    assign twf_m0_real_val[ 47] = 9'sd128; assign twf_m0_imag_val[ 47] = 9'sd0;
    assign twf_m0_real_val[ 48] = 9'sd128; assign twf_m0_imag_val[ 48] = 9'sd0;
    assign twf_m0_real_val[ 49] = 9'sd128; assign twf_m0_imag_val[ 49] = 9'sd0;
    assign twf_m0_real_val[ 50] = 9'sd128; assign twf_m0_imag_val[ 50] = 9'sd0;
    assign twf_m0_real_val[ 51] = 9'sd128; assign twf_m0_imag_val[ 51] = 9'sd0;
    assign twf_m0_real_val[ 52] = 9'sd128; assign twf_m0_imag_val[ 52] = 9'sd0;
    assign twf_m0_real_val[ 53] = 9'sd128; assign twf_m0_imag_val[ 53] = 9'sd0;
    assign twf_m0_real_val[ 54] = 9'sd128; assign twf_m0_imag_val[ 54] = 9'sd0;
    assign twf_m0_real_val[ 55] = 9'sd128; assign twf_m0_imag_val[ 55] = 9'sd0;
    assign twf_m0_real_val[ 56] = 9'sd128; assign twf_m0_imag_val[ 56] = 9'sd0;
    assign twf_m0_real_val[ 57] = 9'sd128; assign twf_m0_imag_val[ 57] = 9'sd0;
    assign twf_m0_real_val[ 58] = 9'sd128; assign twf_m0_imag_val[ 58] = 9'sd0;
    assign twf_m0_real_val[ 59] = 9'sd128; assign twf_m0_imag_val[ 59] = 9'sd0;
    assign twf_m0_real_val[ 60] = 9'sd128; assign twf_m0_imag_val[ 60] = 9'sd0;
    assign twf_m0_real_val[ 61] = 9'sd128; assign twf_m0_imag_val[ 61] = 9'sd0;
    assign twf_m0_real_val[ 62] = 9'sd128; assign twf_m0_imag_val[ 62] = 9'sd0;
    assign twf_m0_real_val[ 63] = 9'sd128; assign twf_m0_imag_val[ 63] = 9'sd0;

    // K3(2) = 4, for nn = 1~64 (index 65~128)
    assign twf_m0_real_val[ 64] = 9'sd128; assign twf_m0_imag_val[ 64] = 9'sd0;
    assign twf_m0_real_val[ 65] = 9'sd128; assign twf_m0_imag_val[ 65] = -9'sd6;
    assign twf_m0_real_val[ 66] = 9'sd127; assign twf_m0_imag_val[ 66] = -9'sd13;
    assign twf_m0_real_val[ 67] = 9'sd127; assign twf_m0_imag_val[ 67] = -9'sd19;
    assign twf_m0_real_val[ 68] = 9'sd126; assign twf_m0_imag_val[ 68] = -9'sd25;
    assign twf_m0_real_val[ 69] = 9'sd124; assign twf_m0_imag_val[ 69] = -9'sd31;
    assign twf_m0_real_val[ 70] = 9'sd122; assign twf_m0_imag_val[ 70] = -9'sd37;
    assign twf_m0_real_val[ 71] = 9'sd121; assign twf_m0_imag_val[ 71] = -9'sd43;
    assign twf_m0_real_val[ 72] = 9'sd118; assign twf_m0_imag_val[ 72] = -9'sd49;
    assign twf_m0_real_val[ 73] = 9'sd116; assign twf_m0_imag_val[ 73] = -9'sd55;
    assign twf_m0_real_val[ 74] = 9'sd113; assign twf_m0_imag_val[ 74] = -9'sd60;
    assign twf_m0_real_val[ 75] = 9'sd110; assign twf_m0_imag_val[ 75] = -9'sd66;
    assign twf_m0_real_val[ 76] = 9'sd106; assign twf_m0_imag_val[ 76] = -9'sd71;
    assign twf_m0_real_val[ 77] = 9'sd103; assign twf_m0_imag_val[ 77] = -9'sd76;
    assign twf_m0_real_val[ 78] = 9'sd99; assign twf_m0_imag_val[ 78] = -9'sd81;
    assign twf_m0_real_val[ 79] = 9'sd95; assign twf_m0_imag_val[ 79] = -9'sd86;
    assign twf_m0_real_val[ 80] = 9'sd91; assign twf_m0_imag_val[ 80] = -9'sd91;
    assign twf_m0_real_val[ 81] = 9'sd86; assign twf_m0_imag_val[ 81] = -9'sd95;
    assign twf_m0_real_val[ 82] = 9'sd81; assign twf_m0_imag_val[ 82] = -9'sd99;
    assign twf_m0_real_val[ 83] = 9'sd76; assign twf_m0_imag_val[ 83] = -9'sd103;
    assign twf_m0_real_val[ 84] = 9'sd71; assign twf_m0_imag_val[ 84] = -9'sd106;
    assign twf_m0_real_val[ 85] = 9'sd66; assign twf_m0_imag_val[ 85] = -9'sd110;
    assign twf_m0_real_val[ 86] = 9'sd60; assign twf_m0_imag_val[ 86] = -9'sd113;
    assign twf_m0_real_val[ 87] = 9'sd55; assign twf_m0_imag_val[ 87] = -9'sd116;
    assign twf_m0_real_val[ 88] = 9'sd49; assign twf_m0_imag_val[ 88] = -9'sd118;
    assign twf_m0_real_val[ 89] = 9'sd43; assign twf_m0_imag_val[ 89] = -9'sd121;
    assign twf_m0_real_val[ 90] = 9'sd37; assign twf_m0_imag_val[ 90] = -9'sd122;
    assign twf_m0_real_val[ 91] = 9'sd31; assign twf_m0_imag_val[ 91] = -9'sd124;
    assign twf_m0_real_val[ 92] = 9'sd25; assign twf_m0_imag_val[ 92] = -9'sd126;
    assign twf_m0_real_val[ 93] = 9'sd19; assign twf_m0_imag_val[ 93] = -9'sd127;
    assign twf_m0_real_val[ 94] = 9'sd13; assign twf_m0_imag_val[ 94] = -9'sd127;
    assign twf_m0_real_val[ 95] = 9'sd6; assign twf_m0_imag_val[ 95] = -9'sd128;
    assign twf_m0_real_val[ 96] = 9'sd0; assign twf_m0_imag_val[ 96] = -9'sd128;
    assign twf_m0_real_val[ 97] = -9'sd6; assign twf_m0_imag_val[ 97] = -9'sd128;
    assign twf_m0_real_val[ 98] = -9'sd13; assign twf_m0_imag_val[ 98] = -9'sd127;
    assign twf_m0_real_val[ 99] = -9'sd19; assign twf_m0_imag_val[ 99] = -9'sd127;
    assign twf_m0_real_val[100] = -9'sd25; assign twf_m0_imag_val[100] = -9'sd126;
    assign twf_m0_real_val[101] = -9'sd31; assign twf_m0_imag_val[101] = -9'sd124;
    assign twf_m0_real_val[102] = -9'sd37; assign twf_m0_imag_val[102] = -9'sd122;
    assign twf_m0_real_val[103] = -9'sd43; assign twf_m0_imag_val[103] = -9'sd121;
    assign twf_m0_real_val[104] = -9'sd49; assign twf_m0_imag_val[104] = -9'sd118;
    assign twf_m0_real_val[105] = -9'sd55; assign twf_m0_imag_val[105] = -9'sd116;
    assign twf_m0_real_val[106] = -9'sd60; assign twf_m0_imag_val[106] = -9'sd113;
    assign twf_m0_real_val[107] = -9'sd66; assign twf_m0_imag_val[107] = -9'sd110;
    assign twf_m0_real_val[108] = -9'sd71; assign twf_m0_imag_val[108] = -9'sd106;
    assign twf_m0_real_val[109] = -9'sd76; assign twf_m0_imag_val[109] = -9'sd103;
    assign twf_m0_real_val[110] = -9'sd81; assign twf_m0_imag_val[110] = -9'sd99;
    assign twf_m0_real_val[111] = -9'sd86; assign twf_m0_imag_val[111] = -9'sd95;
    assign twf_m0_real_val[112] = -9'sd91; assign twf_m0_imag_val[112] = -9'sd91;
    assign twf_m0_real_val[113] = -9'sd95; assign twf_m0_imag_val[113] = -9'sd86;
    assign twf_m0_real_val[114] = -9'sd99; assign twf_m0_imag_val[114] = -9'sd81;
    assign twf_m0_real_val[115] = -9'sd103; assign twf_m0_imag_val[115] = -9'sd76;
    assign twf_m0_real_val[116] = -9'sd106; assign twf_m0_imag_val[116] = -9'sd71;
    assign twf_m0_real_val[117] = -9'sd110; assign twf_m0_imag_val[117] = -9'sd66;
    assign twf_m0_real_val[118] = -9'sd113; assign twf_m0_imag_val[118] = -9'sd60;
    assign twf_m0_real_val[119] = -9'sd116; assign twf_m0_imag_val[119] = -9'sd55;
    assign twf_m0_real_val[120] = -9'sd118; assign twf_m0_imag_val[120] = -9'sd49;
    assign twf_m0_real_val[121] = -9'sd121; assign twf_m0_imag_val[121] = -9'sd43;
    assign twf_m0_real_val[122] = -9'sd122; assign twf_m0_imag_val[122] = -9'sd37;
    assign twf_m0_real_val[123] = -9'sd124; assign twf_m0_imag_val[123] = -9'sd31;
    assign twf_m0_real_val[124] = -9'sd126; assign twf_m0_imag_val[124] = -9'sd25;
    assign twf_m0_real_val[125] = -9'sd127; assign twf_m0_imag_val[125] = -9'sd19;
    assign twf_m0_real_val[126] = -9'sd127; assign twf_m0_imag_val[126] = -9'sd13;
    assign twf_m0_real_val[127] = -9'sd128; assign twf_m0_imag_val[127] = -9'sd6;

    // K3(3) = 2, for nn = 1~64 (index 129~192)
    assign twf_m0_real_val[128] = 9'sd128; assign twf_m0_imag_val[128] = 9'sd0;
    assign twf_m0_real_val[129] = 9'sd128; assign twf_m0_imag_val[129] = -9'sd3;
    assign twf_m0_real_val[130] = 9'sd128; assign twf_m0_imag_val[130] = -9'sd6;
    assign twf_m0_real_val[131] = 9'sd128; assign twf_m0_imag_val[131] = -9'sd9;
    assign twf_m0_real_val[132] = 9'sd127; assign twf_m0_imag_val[132] = -9'sd13;
    assign twf_m0_real_val[133] = 9'sd127; assign twf_m0_imag_val[133] = -9'sd16;
    assign twf_m0_real_val[134] = 9'sd127; assign twf_m0_imag_val[134] = -9'sd19;
    assign twf_m0_real_val[135] = 9'sd126; assign twf_m0_imag_val[135] = -9'sd22;
    assign twf_m0_real_val[136] = 9'sd126; assign twf_m0_imag_val[136] = -9'sd25;
    assign twf_m0_real_val[137] = 9'sd125; assign twf_m0_imag_val[137] = -9'sd28;
    assign twf_m0_real_val[138] = 9'sd124; assign twf_m0_imag_val[138] = -9'sd31;
    assign twf_m0_real_val[139] = 9'sd123; assign twf_m0_imag_val[139] = -9'sd34;
    assign twf_m0_real_val[140] = 9'sd122; assign twf_m0_imag_val[140] = -9'sd37;
    assign twf_m0_real_val[141] = 9'sd122; assign twf_m0_imag_val[141] = -9'sd40;
    assign twf_m0_real_val[142] = 9'sd121; assign twf_m0_imag_val[142] = -9'sd43;
    assign twf_m0_real_val[143] = 9'sd119; assign twf_m0_imag_val[143] = -9'sd46;
    assign twf_m0_real_val[144] = 9'sd118; assign twf_m0_imag_val[144] = -9'sd49;
    assign twf_m0_real_val[145] = 9'sd117; assign twf_m0_imag_val[145] = -9'sd52;
    assign twf_m0_real_val[146] = 9'sd116; assign twf_m0_imag_val[146] = -9'sd55;
    assign twf_m0_real_val[147] = 9'sd114; assign twf_m0_imag_val[147] = -9'sd58;
    assign twf_m0_real_val[148] = 9'sd113; assign twf_m0_imag_val[148] = -9'sd60;
    assign twf_m0_real_val[149] = 9'sd111; assign twf_m0_imag_val[149] = -9'sd63;
    assign twf_m0_real_val[150] = 9'sd110; assign twf_m0_imag_val[150] = -9'sd66;
    assign twf_m0_real_val[151] = 9'sd108; assign twf_m0_imag_val[151] = -9'sd68;
    assign twf_m0_real_val[152] = 9'sd106; assign twf_m0_imag_val[152] = -9'sd71;
    assign twf_m0_real_val[153] = 9'sd105; assign twf_m0_imag_val[153] = -9'sd74;
    assign twf_m0_real_val[154] = 9'sd103; assign twf_m0_imag_val[154] = -9'sd76;
    assign twf_m0_real_val[155] = 9'sd101; assign twf_m0_imag_val[155] = -9'sd79;
    assign twf_m0_real_val[156] = 9'sd99; assign twf_m0_imag_val[156] = -9'sd81;
    assign twf_m0_real_val[157] = 9'sd97; assign twf_m0_imag_val[157] = -9'sd84;
    assign twf_m0_real_val[158] = 9'sd95; assign twf_m0_imag_val[158] = -9'sd86;
    assign twf_m0_real_val[159] = 9'sd93; assign twf_m0_imag_val[159] = -9'sd88;
    assign twf_m0_real_val[160] = 9'sd91; assign twf_m0_imag_val[160] = -9'sd91;
    assign twf_m0_real_val[161] = 9'sd88; assign twf_m0_imag_val[161] = -9'sd93;
    assign twf_m0_real_val[162] = 9'sd86; assign twf_m0_imag_val[162] = -9'sd95;
    assign twf_m0_real_val[163] = 9'sd84; assign twf_m0_imag_val[163] = -9'sd97;
    assign twf_m0_real_val[164] = 9'sd81; assign twf_m0_imag_val[164] = -9'sd99;
    assign twf_m0_real_val[165] = 9'sd79; assign twf_m0_imag_val[165] = -9'sd101;
    assign twf_m0_real_val[166] = 9'sd76; assign twf_m0_imag_val[166] = -9'sd103;
    assign twf_m0_real_val[167] = 9'sd74; assign twf_m0_imag_val[167] = -9'sd105;
    assign twf_m0_real_val[168] = 9'sd71; assign twf_m0_imag_val[168] = -9'sd106;
    assign twf_m0_real_val[169] = 9'sd68; assign twf_m0_imag_val[169] = -9'sd108;
    assign twf_m0_real_val[170] = 9'sd66; assign twf_m0_imag_val[170] = -9'sd110;
    assign twf_m0_real_val[171] = 9'sd63; assign twf_m0_imag_val[171] = -9'sd111;
    assign twf_m0_real_val[172] = 9'sd60; assign twf_m0_imag_val[172] = -9'sd113;
    assign twf_m0_real_val[173] = 9'sd58; assign twf_m0_imag_val[173] = -9'sd114;
    assign twf_m0_real_val[174] = 9'sd55; assign twf_m0_imag_val[174] = -9'sd116;
    assign twf_m0_real_val[175] = 9'sd52; assign twf_m0_imag_val[175] = -9'sd117;
    assign twf_m0_real_val[176] = 9'sd49; assign twf_m0_imag_val[176] = -9'sd118;
    assign twf_m0_real_val[177] = 9'sd46; assign twf_m0_imag_val[177] = -9'sd119;
    assign twf_m0_real_val[178] = 9'sd43; assign twf_m0_imag_val[178] = -9'sd121;
    assign twf_m0_real_val[179] = 9'sd40; assign twf_m0_imag_val[179] = -9'sd122;
    assign twf_m0_real_val[180] = 9'sd37; assign twf_m0_imag_val[180] = -9'sd122;
    assign twf_m0_real_val[181] = 9'sd34; assign twf_m0_imag_val[181] = -9'sd123;
    assign twf_m0_real_val[182] = 9'sd31; assign twf_m0_imag_val[182] = -9'sd124;
    assign twf_m0_real_val[183] = 9'sd28; assign twf_m0_imag_val[183] = -9'sd125;
    assign twf_m0_real_val[184] = 9'sd25; assign twf_m0_imag_val[184] = -9'sd126;
    assign twf_m0_real_val[185] = 9'sd22; assign twf_m0_imag_val[185] = -9'sd126;
    assign twf_m0_real_val[186] = 9'sd19; assign twf_m0_imag_val[186] = -9'sd127;
    assign twf_m0_real_val[187] = 9'sd16; assign twf_m0_imag_val[187] = -9'sd127;
    assign twf_m0_real_val[188] = 9'sd13; assign twf_m0_imag_val[188] = -9'sd127;
    assign twf_m0_real_val[189] = 9'sd9; assign twf_m0_imag_val[189] = -9'sd128;
    assign twf_m0_real_val[190] = 9'sd6; assign twf_m0_imag_val[190] = -9'sd128;
    assign twf_m0_real_val[191] = 9'sd3; assign twf_m0_imag_val[191] = -9'sd128;

    // K3(4) = 6, for nn = 1~64 (index 193~256)
    assign twf_m0_real_val[192] = 9'sd128; assign twf_m0_imag_val[192] = 9'sd0;
    assign twf_m0_real_val[193] = 9'sd128; assign twf_m0_imag_val[193] = -9'sd9;
    assign twf_m0_real_val[194] = 9'sd127; assign twf_m0_imag_val[194] = -9'sd19;
    assign twf_m0_real_val[195] = 9'sd125; assign twf_m0_imag_val[195] = -9'sd28;
    assign twf_m0_real_val[196] = 9'sd122; assign twf_m0_imag_val[196] = -9'sd37;
    assign twf_m0_real_val[197] = 9'sd119; assign twf_m0_imag_val[197] = -9'sd46;
    assign twf_m0_real_val[198] = 9'sd116; assign twf_m0_imag_val[198] = -9'sd55;
    assign twf_m0_real_val[199] = 9'sd111; assign twf_m0_imag_val[199] = -9'sd63;
    assign twf_m0_real_val[200] = 9'sd106; assign twf_m0_imag_val[200] = -9'sd71;
    assign twf_m0_real_val[201] = 9'sd101; assign twf_m0_imag_val[201] = -9'sd79;
    assign twf_m0_real_val[202] = 9'sd95; assign twf_m0_imag_val[202] = -9'sd86;
    assign twf_m0_real_val[203] = 9'sd88; assign twf_m0_imag_val[203] = -9'sd93;
    assign twf_m0_real_val[204] = 9'sd81; assign twf_m0_imag_val[204] = -9'sd99;
    assign twf_m0_real_val[205] = 9'sd74; assign twf_m0_imag_val[205] = -9'sd105;
    assign twf_m0_real_val[206] = 9'sd66; assign twf_m0_imag_val[206] = -9'sd110;
    assign twf_m0_real_val[207] = 9'sd58; assign twf_m0_imag_val[207] = -9'sd114;
    assign twf_m0_real_val[208] = 9'sd49; assign twf_m0_imag_val[208] = -9'sd118;
    assign twf_m0_real_val[209] = 9'sd40; assign twf_m0_imag_val[209] = -9'sd122;
    assign twf_m0_real_val[210] = 9'sd31; assign twf_m0_imag_val[210] = -9'sd124;
    assign twf_m0_real_val[211] = 9'sd22; assign twf_m0_imag_val[211] = -9'sd126;
    assign twf_m0_real_val[212] = 9'sd13; assign twf_m0_imag_val[212] = -9'sd127;
    assign twf_m0_real_val[213] = 9'sd3; assign twf_m0_imag_val[213] = -9'sd128;
    assign twf_m0_real_val[214] = -9'sd6; assign twf_m0_imag_val[214] = -9'sd128;
    assign twf_m0_real_val[215] = -9'sd16; assign twf_m0_imag_val[215] = -9'sd127;
    assign twf_m0_real_val[216] = -9'sd25; assign twf_m0_imag_val[216] = -9'sd126;
    assign twf_m0_real_val[217] = -9'sd34; assign twf_m0_imag_val[217] = -9'sd123;
    assign twf_m0_real_val[218] = -9'sd43; assign twf_m0_imag_val[218] = -9'sd121;
    assign twf_m0_real_val[219] = -9'sd52; assign twf_m0_imag_val[219] = -9'sd117;
    assign twf_m0_real_val[220] = -9'sd60; assign twf_m0_imag_val[220] = -9'sd113;
    assign twf_m0_real_val[221] = -9'sd68; assign twf_m0_imag_val[221] = -9'sd108;
    assign twf_m0_real_val[222] = -9'sd76; assign twf_m0_imag_val[222] = -9'sd103;
    assign twf_m0_real_val[223] = -9'sd84; assign twf_m0_imag_val[223] = -9'sd97;
    assign twf_m0_real_val[224] = -9'sd91; assign twf_m0_imag_val[224] = -9'sd91;
    assign twf_m0_real_val[225] = -9'sd97; assign twf_m0_imag_val[225] = -9'sd84;
    assign twf_m0_real_val[226] = -9'sd103; assign twf_m0_imag_val[226] = -9'sd76;
    assign twf_m0_real_val[227] = -9'sd108; assign twf_m0_imag_val[227] = -9'sd68;
    assign twf_m0_real_val[228] = -9'sd113; assign twf_m0_imag_val[228] = -9'sd60;
    assign twf_m0_real_val[229] = -9'sd117; assign twf_m0_imag_val[229] = -9'sd52;
    assign twf_m0_real_val[230] = -9'sd121; assign twf_m0_imag_val[230] = -9'sd43;
    assign twf_m0_real_val[231] = -9'sd123; assign twf_m0_imag_val[231] = -9'sd34;
    assign twf_m0_real_val[232] = -9'sd126; assign twf_m0_imag_val[232] = -9'sd25;
    assign twf_m0_real_val[233] = -9'sd127; assign twf_m0_imag_val[233] = -9'sd16;
    assign twf_m0_real_val[234] = -9'sd128; assign twf_m0_imag_val[234] = -9'sd6;
    assign twf_m0_real_val[235] = -9'sd128; assign twf_m0_imag_val[235] = 9'sd3;
    assign twf_m0_real_val[236] = -9'sd127; assign twf_m0_imag_val[236] = 9'sd13;
    assign twf_m0_real_val[237] = -9'sd126; assign twf_m0_imag_val[237] = 9'sd22;
    assign twf_m0_real_val[238] = -9'sd124; assign twf_m0_imag_val[238] = 9'sd31;
    assign twf_m0_real_val[239] = -9'sd122; assign twf_m0_imag_val[239] = 9'sd40;
    assign twf_m0_real_val[240] = -9'sd118; assign twf_m0_imag_val[240] = 9'sd49;
    assign twf_m0_real_val[241] = -9'sd114; assign twf_m0_imag_val[241] = 9'sd58;
    assign twf_m0_real_val[242] = -9'sd110; assign twf_m0_imag_val[242] = 9'sd66;
    assign twf_m0_real_val[243] = -9'sd105; assign twf_m0_imag_val[243] = 9'sd74;
    assign twf_m0_real_val[244] = -9'sd99; assign twf_m0_imag_val[244] = 9'sd81;
    assign twf_m0_real_val[245] = -9'sd93; assign twf_m0_imag_val[245] = 9'sd88;
    assign twf_m0_real_val[246] = -9'sd86; assign twf_m0_imag_val[246] = 9'sd95;
    assign twf_m0_real_val[247] = -9'sd79; assign twf_m0_imag_val[247] = 9'sd101;
    assign twf_m0_real_val[248] = -9'sd71; assign twf_m0_imag_val[248] = 9'sd106;
    assign twf_m0_real_val[249] = -9'sd63; assign twf_m0_imag_val[249] = 9'sd111;
    assign twf_m0_real_val[250] = -9'sd55; assign twf_m0_imag_val[250] = 9'sd116;
    assign twf_m0_real_val[251] = -9'sd46; assign twf_m0_imag_val[251] = 9'sd119;
    assign twf_m0_real_val[252] = -9'sd37; assign twf_m0_imag_val[252] = 9'sd122;
    assign twf_m0_real_val[253] = -9'sd28; assign twf_m0_imag_val[253] = 9'sd125;
    assign twf_m0_real_val[254] = -9'sd19; assign twf_m0_imag_val[254] = 9'sd127;
    assign twf_m0_real_val[255] = -9'sd9; assign twf_m0_imag_val[255] = 9'sd128;

    // K3(5) = 1, for nn = 1~64 (index 257~320)
    assign twf_m0_real_val[256] = 9'sd128; assign twf_m0_imag_val[256] = 9'sd0;
    assign twf_m0_real_val[257] = 9'sd128; assign twf_m0_imag_val[257] = -9'sd2;
    assign twf_m0_real_val[258] = 9'sd128; assign twf_m0_imag_val[258] = -9'sd3;
    assign twf_m0_real_val[259] = 9'sd128; assign twf_m0_imag_val[259] = -9'sd5;
    assign twf_m0_real_val[260] = 9'sd128; assign twf_m0_imag_val[260] = -9'sd6;
    assign twf_m0_real_val[261] = 9'sd128; assign twf_m0_imag_val[261] = -9'sd8;
    assign twf_m0_real_val[262] = 9'sd128; assign twf_m0_imag_val[262] = -9'sd9;
    assign twf_m0_real_val[263] = 9'sd128; assign twf_m0_imag_val[263] = -9'sd11;
    assign twf_m0_real_val[264] = 9'sd127; assign twf_m0_imag_val[264] = -9'sd13;
    assign twf_m0_real_val[265] = 9'sd127; assign twf_m0_imag_val[265] = -9'sd14;
    assign twf_m0_real_val[266] = 9'sd127; assign twf_m0_imag_val[266] = -9'sd16;
    assign twf_m0_real_val[267] = 9'sd127; assign twf_m0_imag_val[267] = -9'sd17;
    assign twf_m0_real_val[268] = 9'sd127; assign twf_m0_imag_val[268] = -9'sd19;
    assign twf_m0_real_val[269] = 9'sd126; assign twf_m0_imag_val[269] = -9'sd20;
    assign twf_m0_real_val[270] = 9'sd126; assign twf_m0_imag_val[270] = -9'sd22;
    assign twf_m0_real_val[271] = 9'sd126; assign twf_m0_imag_val[271] = -9'sd23;
    assign twf_m0_real_val[272] = 9'sd126; assign twf_m0_imag_val[272] = -9'sd25;
    assign twf_m0_real_val[273] = 9'sd125; assign twf_m0_imag_val[273] = -9'sd27;
    assign twf_m0_real_val[274] = 9'sd125; assign twf_m0_imag_val[274] = -9'sd28;
    assign twf_m0_real_val[275] = 9'sd125; assign twf_m0_imag_val[275] = -9'sd30;
    assign twf_m0_real_val[276] = 9'sd124; assign twf_m0_imag_val[276] = -9'sd31;
    assign twf_m0_real_val[277] = 9'sd124; assign twf_m0_imag_val[277] = -9'sd33;
    assign twf_m0_real_val[278] = 9'sd123; assign twf_m0_imag_val[278] = -9'sd34;
    assign twf_m0_real_val[279] = 9'sd123; assign twf_m0_imag_val[279] = -9'sd36;
    assign twf_m0_real_val[280] = 9'sd122; assign twf_m0_imag_val[280] = -9'sd37;
    assign twf_m0_real_val[281] = 9'sd122; assign twf_m0_imag_val[281] = -9'sd39;
    assign twf_m0_real_val[282] = 9'sd122; assign twf_m0_imag_val[282] = -9'sd40;
    assign twf_m0_real_val[283] = 9'sd121; assign twf_m0_imag_val[283] = -9'sd42;
    assign twf_m0_real_val[284] = 9'sd121; assign twf_m0_imag_val[284] = -9'sd43;
    assign twf_m0_real_val[285] = 9'sd120; assign twf_m0_imag_val[285] = -9'sd45;
    assign twf_m0_real_val[286] = 9'sd119; assign twf_m0_imag_val[286] = -9'sd46;
    assign twf_m0_real_val[287] = 9'sd119; assign twf_m0_imag_val[287] = -9'sd48;
    assign twf_m0_real_val[288] = 9'sd118; assign twf_m0_imag_val[288] = -9'sd49;
    assign twf_m0_real_val[289] = 9'sd118; assign twf_m0_imag_val[289] = -9'sd50;
    assign twf_m0_real_val[290] = 9'sd117; assign twf_m0_imag_val[290] = -9'sd52;
    assign twf_m0_real_val[291] = 9'sd116; assign twf_m0_imag_val[291] = -9'sd53;
    assign twf_m0_real_val[292] = 9'sd116; assign twf_m0_imag_val[292] = -9'sd55;
    assign twf_m0_real_val[293] = 9'sd115; assign twf_m0_imag_val[293] = -9'sd56;
    assign twf_m0_real_val[294] = 9'sd114; assign twf_m0_imag_val[294] = -9'sd58;
    assign twf_m0_real_val[295] = 9'sd114; assign twf_m0_imag_val[295] = -9'sd59;
    assign twf_m0_real_val[296] = 9'sd113; assign twf_m0_imag_val[296] = -9'sd60;
    assign twf_m0_real_val[297] = 9'sd112; assign twf_m0_imag_val[297] = -9'sd62;
    assign twf_m0_real_val[298] = 9'sd111; assign twf_m0_imag_val[298] = -9'sd63;
    assign twf_m0_real_val[299] = 9'sd111; assign twf_m0_imag_val[299] = -9'sd64;
    assign twf_m0_real_val[300] = 9'sd110; assign twf_m0_imag_val[300] = -9'sd66;
    assign twf_m0_real_val[301] = 9'sd109; assign twf_m0_imag_val[301] = -9'sd67;
    assign twf_m0_real_val[302] = 9'sd108; assign twf_m0_imag_val[302] = -9'sd68;
    assign twf_m0_real_val[303] = 9'sd107; assign twf_m0_imag_val[303] = -9'sd70;
    assign twf_m0_real_val[304] = 9'sd106; assign twf_m0_imag_val[304] = -9'sd71;
    assign twf_m0_real_val[305] = 9'sd106; assign twf_m0_imag_val[305] = -9'sd72;
    assign twf_m0_real_val[306] = 9'sd105; assign twf_m0_imag_val[306] = -9'sd74;
    assign twf_m0_real_val[307] = 9'sd104; assign twf_m0_imag_val[307] = -9'sd75;
    assign twf_m0_real_val[308] = 9'sd103; assign twf_m0_imag_val[308] = -9'sd76;
    assign twf_m0_real_val[309] = 9'sd102; assign twf_m0_imag_val[309] = -9'sd78;
    assign twf_m0_real_val[310] = 9'sd101; assign twf_m0_imag_val[310] = -9'sd79;
    assign twf_m0_real_val[311] = 9'sd100; assign twf_m0_imag_val[311] = -9'sd80;
    assign twf_m0_real_val[312] = 9'sd99; assign twf_m0_imag_val[312] = -9'sd81;
    assign twf_m0_real_val[313] = 9'sd98; assign twf_m0_imag_val[313] = -9'sd82;
    assign twf_m0_real_val[314] = 9'sd97; assign twf_m0_imag_val[314] = -9'sd84;
    assign twf_m0_real_val[315] = 9'sd96; assign twf_m0_imag_val[315] = -9'sd85;
    assign twf_m0_real_val[316] = 9'sd95; assign twf_m0_imag_val[316] = -9'sd86;
    assign twf_m0_real_val[317] = 9'sd94; assign twf_m0_imag_val[317] = -9'sd87;
    assign twf_m0_real_val[318] = 9'sd93; assign twf_m0_imag_val[318] = -9'sd88;
    assign twf_m0_real_val[319] = 9'sd92; assign twf_m0_imag_val[319] = -9'sd89;

    // K3(6) = 5, for nn = 1~64 (index 321~384)
    assign twf_m0_real_val[320] = 9'sd128; assign twf_m0_imag_val[320] = 9'sd0;
    assign twf_m0_real_val[321] = 9'sd128; assign twf_m0_imag_val[321] = -9'sd8;
    assign twf_m0_real_val[322] = 9'sd127; assign twf_m0_imag_val[322] = -9'sd16;
    assign twf_m0_real_val[323] = 9'sd126; assign twf_m0_imag_val[323] = -9'sd23;
    assign twf_m0_real_val[324] = 9'sd124; assign twf_m0_imag_val[324] = -9'sd31;
    assign twf_m0_real_val[325] = 9'sd122; assign twf_m0_imag_val[325] = -9'sd39;
    assign twf_m0_real_val[326] = 9'sd119; assign twf_m0_imag_val[326] = -9'sd46;
    assign twf_m0_real_val[327] = 9'sd116; assign twf_m0_imag_val[327] = -9'sd53;
    assign twf_m0_real_val[328] = 9'sd113; assign twf_m0_imag_val[328] = -9'sd60;
    assign twf_m0_real_val[329] = 9'sd109; assign twf_m0_imag_val[329] = -9'sd67;
    assign twf_m0_real_val[330] = 9'sd105; assign twf_m0_imag_val[330] = -9'sd74;
    assign twf_m0_real_val[331] = 9'sd100; assign twf_m0_imag_val[331] = -9'sd80;
    assign twf_m0_real_val[332] = 9'sd95; assign twf_m0_imag_val[332] = -9'sd86;
    assign twf_m0_real_val[333] = 9'sd89; assign twf_m0_imag_val[333] = -9'sd92;
    assign twf_m0_real_val[334] = 9'sd84; assign twf_m0_imag_val[334] = -9'sd97;
    assign twf_m0_real_val[335] = 9'sd78; assign twf_m0_imag_val[335] = -9'sd102;
    assign twf_m0_real_val[336] = 9'sd71; assign twf_m0_imag_val[336] = -9'sd106;
    assign twf_m0_real_val[337] = 9'sd64; assign twf_m0_imag_val[337] = -9'sd111;
    assign twf_m0_real_val[338] = 9'sd58; assign twf_m0_imag_val[338] = -9'sd114;
    assign twf_m0_real_val[339] = 9'sd50; assign twf_m0_imag_val[339] = -9'sd118;
    assign twf_m0_real_val[340] = 9'sd43; assign twf_m0_imag_val[340] = -9'sd121;
    assign twf_m0_real_val[341] = 9'sd36; assign twf_m0_imag_val[341] = -9'sd123;
    assign twf_m0_real_val[342] = 9'sd28; assign twf_m0_imag_val[342] = -9'sd125;
    assign twf_m0_real_val[343] = 9'sd20; assign twf_m0_imag_val[343] = -9'sd126;
    assign twf_m0_real_val[344] = 9'sd13; assign twf_m0_imag_val[344] = -9'sd127;
    assign twf_m0_real_val[345] = 9'sd5; assign twf_m0_imag_val[345] = -9'sd128;
    assign twf_m0_real_val[346] = -9'sd3; assign twf_m0_imag_val[346] = -9'sd128;
    assign twf_m0_real_val[347] = -9'sd11; assign twf_m0_imag_val[347] = -9'sd128;
    assign twf_m0_real_val[348] = -9'sd19; assign twf_m0_imag_val[348] = -9'sd127;
    assign twf_m0_real_val[349] = -9'sd27; assign twf_m0_imag_val[349] = -9'sd125;
    assign twf_m0_real_val[350] = -9'sd34; assign twf_m0_imag_val[350] = -9'sd123;
    assign twf_m0_real_val[351] = -9'sd42; assign twf_m0_imag_val[351] = -9'sd121;
    assign twf_m0_real_val[352] = -9'sd49; assign twf_m0_imag_val[352] = -9'sd118;
    assign twf_m0_real_val[353] = -9'sd56; assign twf_m0_imag_val[353] = -9'sd115;
    assign twf_m0_real_val[354] = -9'sd63; assign twf_m0_imag_val[354] = -9'sd111;
    assign twf_m0_real_val[355] = -9'sd70; assign twf_m0_imag_val[355] = -9'sd107;
    assign twf_m0_real_val[356] = -9'sd76; assign twf_m0_imag_val[356] = -9'sd103;
    assign twf_m0_real_val[357] = -9'sd82; assign twf_m0_imag_val[357] = -9'sd98;
    assign twf_m0_real_val[358] = -9'sd88; assign twf_m0_imag_val[358] = -9'sd93;
    assign twf_m0_real_val[359] = -9'sd94; assign twf_m0_imag_val[359] = -9'sd87;
    assign twf_m0_real_val[360] = -9'sd99; assign twf_m0_imag_val[360] = -9'sd81;
    assign twf_m0_real_val[361] = -9'sd104; assign twf_m0_imag_val[361] = -9'sd75;
    assign twf_m0_real_val[362] = -9'sd108; assign twf_m0_imag_val[362] = -9'sd68;
    assign twf_m0_real_val[363] = -9'sd112; assign twf_m0_imag_val[363] = -9'sd62;
    assign twf_m0_real_val[364] = -9'sd116; assign twf_m0_imag_val[364] = -9'sd55;
    assign twf_m0_real_val[365] = -9'sd119; assign twf_m0_imag_val[365] = -9'sd48;
    assign twf_m0_real_val[366] = -9'sd122; assign twf_m0_imag_val[366] = -9'sd40;
    assign twf_m0_real_val[367] = -9'sd124; assign twf_m0_imag_val[367] = -9'sd33;
    assign twf_m0_real_val[368] = -9'sd126; assign twf_m0_imag_val[368] = -9'sd25;
    assign twf_m0_real_val[369] = -9'sd127; assign twf_m0_imag_val[369] = -9'sd17;
    assign twf_m0_real_val[370] = -9'sd128; assign twf_m0_imag_val[370] = -9'sd9;
    assign twf_m0_real_val[371] = -9'sd128; assign twf_m0_imag_val[371] = -9'sd2;
    assign twf_m0_real_val[372] = -9'sd128; assign twf_m0_imag_val[372] = 9'sd6;
    assign twf_m0_real_val[373] = -9'sd127; assign twf_m0_imag_val[373] = 9'sd14;
    assign twf_m0_real_val[374] = -9'sd126; assign twf_m0_imag_val[374] = 9'sd22;
    assign twf_m0_real_val[375] = -9'sd125; assign twf_m0_imag_val[375] = 9'sd30;
    assign twf_m0_real_val[376] = -9'sd122; assign twf_m0_imag_val[376] = 9'sd37;
    assign twf_m0_real_val[377] = -9'sd120; assign twf_m0_imag_val[377] = 9'sd45;
    assign twf_m0_real_val[378] = -9'sd117; assign twf_m0_imag_val[378] = 9'sd52;
    assign twf_m0_real_val[379] = -9'sd114; assign twf_m0_imag_val[379] = 9'sd59;
    assign twf_m0_real_val[380] = -9'sd110; assign twf_m0_imag_val[380] = 9'sd66;
    assign twf_m0_real_val[381] = -9'sd106; assign twf_m0_imag_val[381] = 9'sd72;
    assign twf_m0_real_val[382] = -9'sd101; assign twf_m0_imag_val[382] = 9'sd79;
    assign twf_m0_real_val[383] = -9'sd96; assign twf_m0_imag_val[383] = 9'sd85;

    // K3(7) = 3, for nn = 1~64 (index 385~448)
    assign twf_m0_real_val[384] = 9'sd128; assign twf_m0_imag_val[384] = 9'sd0;
    assign twf_m0_real_val[385] = 9'sd128; assign twf_m0_imag_val[385] = -9'sd5;
    assign twf_m0_real_val[386] = 9'sd128; assign twf_m0_imag_val[386] = -9'sd9;
    assign twf_m0_real_val[387] = 9'sd127; assign twf_m0_imag_val[387] = -9'sd14;
    assign twf_m0_real_val[388] = 9'sd127; assign twf_m0_imag_val[388] = -9'sd19;
    assign twf_m0_real_val[389] = 9'sd126; assign twf_m0_imag_val[389] = -9'sd23;
    assign twf_m0_real_val[390] = 9'sd125; assign twf_m0_imag_val[390] = -9'sd28;
    assign twf_m0_real_val[391] = 9'sd124; assign twf_m0_imag_val[391] = -9'sd33;
    assign twf_m0_real_val[392] = 9'sd122; assign twf_m0_imag_val[392] = -9'sd37;
    assign twf_m0_real_val[393] = 9'sd121; assign twf_m0_imag_val[393] = -9'sd42;
    assign twf_m0_real_val[394] = 9'sd119; assign twf_m0_imag_val[394] = -9'sd46;
    assign twf_m0_real_val[395] = 9'sd118; assign twf_m0_imag_val[395] = -9'sd50;
    assign twf_m0_real_val[396] = 9'sd116; assign twf_m0_imag_val[396] = -9'sd55;
    assign twf_m0_real_val[397] = 9'sd114; assign twf_m0_imag_val[397] = -9'sd59;
    assign twf_m0_real_val[398] = 9'sd111; assign twf_m0_imag_val[398] = -9'sd63;
    assign twf_m0_real_val[399] = 9'sd109; assign twf_m0_imag_val[399] = -9'sd67;
    assign twf_m0_real_val[400] = 9'sd106; assign twf_m0_imag_val[400] = -9'sd71;
    assign twf_m0_real_val[401] = 9'sd104; assign twf_m0_imag_val[401] = -9'sd75;
    assign twf_m0_real_val[402] = 9'sd101; assign twf_m0_imag_val[402] = -9'sd79;
    assign twf_m0_real_val[403] = 9'sd98; assign twf_m0_imag_val[403] = -9'sd82;
    assign twf_m0_real_val[404] = 9'sd95; assign twf_m0_imag_val[404] = -9'sd86;
    assign twf_m0_real_val[405] = 9'sd92; assign twf_m0_imag_val[405] = -9'sd89;
    assign twf_m0_real_val[406] = 9'sd88; assign twf_m0_imag_val[406] = -9'sd93;
    assign twf_m0_real_val[407] = 9'sd85; assign twf_m0_imag_val[407] = -9'sd96;
    assign twf_m0_real_val[408] = 9'sd81; assign twf_m0_imag_val[408] = -9'sd99;
    assign twf_m0_real_val[409] = 9'sd78; assign twf_m0_imag_val[409] = -9'sd102;
    assign twf_m0_real_val[410] = 9'sd74; assign twf_m0_imag_val[410] = -9'sd105;
    assign twf_m0_real_val[411] = 9'sd70; assign twf_m0_imag_val[411] = -9'sd107;
    assign twf_m0_real_val[412] = 9'sd66; assign twf_m0_imag_val[412] = -9'sd110;
    assign twf_m0_real_val[413] = 9'sd62; assign twf_m0_imag_val[413] = -9'sd112;
    assign twf_m0_real_val[414] = 9'sd58; assign twf_m0_imag_val[414] = -9'sd114;
    assign twf_m0_real_val[415] = 9'sd53; assign twf_m0_imag_val[415] = -9'sd116;
    assign twf_m0_real_val[416] = 9'sd49; assign twf_m0_imag_val[416] = -9'sd118;
    assign twf_m0_real_val[417] = 9'sd45; assign twf_m0_imag_val[417] = -9'sd120;
    assign twf_m0_real_val[418] = 9'sd40; assign twf_m0_imag_val[418] = -9'sd122;
    assign twf_m0_real_val[419] = 9'sd36; assign twf_m0_imag_val[419] = -9'sd123;
    assign twf_m0_real_val[420] = 9'sd31; assign twf_m0_imag_val[420] = -9'sd124;
    assign twf_m0_real_val[421] = 9'sd27; assign twf_m0_imag_val[421] = -9'sd125;
    assign twf_m0_real_val[422] = 9'sd22; assign twf_m0_imag_val[422] = -9'sd126;
    assign twf_m0_real_val[423] = 9'sd17; assign twf_m0_imag_val[423] = -9'sd127;
    assign twf_m0_real_val[424] = 9'sd13; assign twf_m0_imag_val[424] = -9'sd127;
    assign twf_m0_real_val[425] = 9'sd8; assign twf_m0_imag_val[425] = -9'sd128;
    assign twf_m0_real_val[426] = 9'sd3; assign twf_m0_imag_val[426] = -9'sd128;
    assign twf_m0_real_val[427] = -9'sd2; assign twf_m0_imag_val[427] = -9'sd128;
    assign twf_m0_real_val[428] = -9'sd6; assign twf_m0_imag_val[428] = -9'sd128;
    assign twf_m0_real_val[429] = -9'sd11; assign twf_m0_imag_val[429] = -9'sd128;
    assign twf_m0_real_val[430] = -9'sd16; assign twf_m0_imag_val[430] = -9'sd127;
    assign twf_m0_real_val[431] = -9'sd20; assign twf_m0_imag_val[431] = -9'sd126;
    assign twf_m0_real_val[432] = -9'sd25; assign twf_m0_imag_val[432] = -9'sd126;
    assign twf_m0_real_val[433] = -9'sd30; assign twf_m0_imag_val[433] = -9'sd125;
    assign twf_m0_real_val[434] = -9'sd34; assign twf_m0_imag_val[434] = -9'sd123;
    assign twf_m0_real_val[435] = -9'sd39; assign twf_m0_imag_val[435] = -9'sd122;
    assign twf_m0_real_val[436] = -9'sd43; assign twf_m0_imag_val[436] = -9'sd121;
    assign twf_m0_real_val[437] = -9'sd48; assign twf_m0_imag_val[437] = -9'sd119;
    assign twf_m0_real_val[438] = -9'sd52; assign twf_m0_imag_val[438] = -9'sd117;
    assign twf_m0_real_val[439] = -9'sd56; assign twf_m0_imag_val[439] = -9'sd115;
    assign twf_m0_real_val[440] = -9'sd60; assign twf_m0_imag_val[440] = -9'sd113;
    assign twf_m0_real_val[441] = -9'sd64; assign twf_m0_imag_val[441] = -9'sd111;
    assign twf_m0_real_val[442] = -9'sd68; assign twf_m0_imag_val[442] = -9'sd108;
    assign twf_m0_real_val[443] = -9'sd72; assign twf_m0_imag_val[443] = -9'sd106;
    assign twf_m0_real_val[444] = -9'sd76; assign twf_m0_imag_val[444] = -9'sd103;
    assign twf_m0_real_val[445] = -9'sd80; assign twf_m0_imag_val[445] = -9'sd100;
    assign twf_m0_real_val[446] = -9'sd84; assign twf_m0_imag_val[446] = -9'sd97;
    assign twf_m0_real_val[447] = -9'sd87; assign twf_m0_imag_val[447] = -9'sd94;

    // K3(8) = 7, for nn = 1~64 (index 449~512)
    assign twf_m0_real_val[448] = 9'sd128; assign twf_m0_imag_val[448] = 9'sd0;
    assign twf_m0_real_val[449] = 9'sd128; assign twf_m0_imag_val[449] = -9'sd11;
    assign twf_m0_real_val[450] = 9'sd126; assign twf_m0_imag_val[450] = -9'sd22;
    assign twf_m0_real_val[451] = 9'sd124; assign twf_m0_imag_val[451] = -9'sd33;
    assign twf_m0_real_val[452] = 9'sd121; assign twf_m0_imag_val[452] = -9'sd43;
    assign twf_m0_real_val[453] = 9'sd116; assign twf_m0_imag_val[453] = -9'sd53;
    assign twf_m0_real_val[454] = 9'sd111; assign twf_m0_imag_val[454] = -9'sd63;
    assign twf_m0_real_val[455] = 9'sd106; assign twf_m0_imag_val[455] = -9'sd72;
    assign twf_m0_real_val[456] = 9'sd99; assign twf_m0_imag_val[456] = -9'sd81;
    assign twf_m0_real_val[457] = 9'sd92; assign twf_m0_imag_val[457] = -9'sd89;
    assign twf_m0_real_val[458] = 9'sd84; assign twf_m0_imag_val[458] = -9'sd97;
    assign twf_m0_real_val[459] = 9'sd75; assign twf_m0_imag_val[459] = -9'sd104;
    assign twf_m0_real_val[460] = 9'sd66; assign twf_m0_imag_val[460] = -9'sd110;
    assign twf_m0_real_val[461] = 9'sd56; assign twf_m0_imag_val[461] = -9'sd115;
    assign twf_m0_real_val[462] = 9'sd46; assign twf_m0_imag_val[462] = -9'sd119;
    assign twf_m0_real_val[463] = 9'sd36; assign twf_m0_imag_val[463] = -9'sd123;
    assign twf_m0_real_val[464] = 9'sd25; assign twf_m0_imag_val[464] = -9'sd126;
    assign twf_m0_real_val[465] = 9'sd14; assign twf_m0_imag_val[465] = -9'sd127;
    assign twf_m0_real_val[466] = 9'sd3; assign twf_m0_imag_val[466] = -9'sd128;
    assign twf_m0_real_val[467] = -9'sd8; assign twf_m0_imag_val[467] = -9'sd128;
    assign twf_m0_real_val[468] = -9'sd19; assign twf_m0_imag_val[468] = -9'sd127;
    assign twf_m0_real_val[469] = -9'sd30; assign twf_m0_imag_val[469] = -9'sd125;
    assign twf_m0_real_val[470] = -9'sd40; assign twf_m0_imag_val[470] = -9'sd122;
    assign twf_m0_real_val[471] = -9'sd50; assign twf_m0_imag_val[471] = -9'sd118;
    assign twf_m0_real_val[472] = -9'sd60; assign twf_m0_imag_val[472] = -9'sd113;
    assign twf_m0_real_val[473] = -9'sd70; assign twf_m0_imag_val[473] = -9'sd107;
    assign twf_m0_real_val[474] = -9'sd79; assign twf_m0_imag_val[474] = -9'sd101;
    assign twf_m0_real_val[475] = -9'sd87; assign twf_m0_imag_val[475] = -9'sd94;
    assign twf_m0_real_val[476] = -9'sd95; assign twf_m0_imag_val[476] = -9'sd86;
    assign twf_m0_real_val[477] = -9'sd102; assign twf_m0_imag_val[477] = -9'sd78;
    assign twf_m0_real_val[478] = -9'sd108; assign twf_m0_imag_val[478] = -9'sd68;
    assign twf_m0_real_val[479] = -9'sd114; assign twf_m0_imag_val[479] = -9'sd59;
    assign twf_m0_real_val[480] = -9'sd118; assign twf_m0_imag_val[480] = -9'sd49;
    assign twf_m0_real_val[481] = -9'sd122; assign twf_m0_imag_val[481] = -9'sd39;
    assign twf_m0_real_val[482] = -9'sd125; assign twf_m0_imag_val[482] = -9'sd28;
    assign twf_m0_real_val[483] = -9'sd127; assign twf_m0_imag_val[483] = -9'sd17;
    assign twf_m0_real_val[484] = -9'sd128; assign twf_m0_imag_val[484] = -9'sd6;
    assign twf_m0_real_val[485] = -9'sd128; assign twf_m0_imag_val[485] = 9'sd5;
    assign twf_m0_real_val[486] = -9'sd127; assign twf_m0_imag_val[486] = 9'sd16;
    assign twf_m0_real_val[487] = -9'sd125; assign twf_m0_imag_val[487] = 9'sd27;
    assign twf_m0_real_val[488] = -9'sd122; assign twf_m0_imag_val[488] = 9'sd37;
    assign twf_m0_real_val[489] = -9'sd119; assign twf_m0_imag_val[489] = 9'sd48;
    assign twf_m0_real_val[490] = -9'sd114; assign twf_m0_imag_val[490] = 9'sd58;
    assign twf_m0_real_val[491] = -9'sd109; assign twf_m0_imag_val[491] = 9'sd67;
    assign twf_m0_real_val[492] = -9'sd103; assign twf_m0_imag_val[492] = 9'sd76;
    assign twf_m0_real_val[493] = -9'sd96; assign twf_m0_imag_val[493] = 9'sd85;
    assign twf_m0_real_val[494] = -9'sd88; assign twf_m0_imag_val[494] = 9'sd93;
    assign twf_m0_real_val[495] = -9'sd80; assign twf_m0_imag_val[495] = 9'sd100;
    assign twf_m0_real_val[496] = -9'sd71; assign twf_m0_imag_val[496] = 9'sd106;
    assign twf_m0_real_val[497] = -9'sd62; assign twf_m0_imag_val[497] = 9'sd112;
    assign twf_m0_real_val[498] = -9'sd52; assign twf_m0_imag_val[498] = 9'sd117;
    assign twf_m0_real_val[499] = -9'sd42; assign twf_m0_imag_val[499] = 9'sd121;
    assign twf_m0_real_val[500] = -9'sd31; assign twf_m0_imag_val[500] = 9'sd124;
    assign twf_m0_real_val[501] = -9'sd20; assign twf_m0_imag_val[501] = 9'sd126;
    assign twf_m0_real_val[502] = -9'sd9; assign twf_m0_imag_val[502] = 9'sd128;
    assign twf_m0_real_val[503] = 9'sd2; assign twf_m0_imag_val[503] = 9'sd128;
    assign twf_m0_real_val[504] = 9'sd13; assign twf_m0_imag_val[504] = 9'sd127;
    assign twf_m0_real_val[505] = 9'sd23; assign twf_m0_imag_val[505] = 9'sd126;
    assign twf_m0_real_val[506] = 9'sd34; assign twf_m0_imag_val[506] = 9'sd123;
    assign twf_m0_real_val[507] = 9'sd45; assign twf_m0_imag_val[507] = 9'sd120;
    assign twf_m0_real_val[508] = 9'sd55; assign twf_m0_imag_val[508] = 9'sd116;
    assign twf_m0_real_val[509] = 9'sd64; assign twf_m0_imag_val[509] = 9'sd111;
    assign twf_m0_real_val[510] = 9'sd74; assign twf_m0_imag_val[510] = 9'sd105;
    assign twf_m0_real_val[511] = 9'sd82; assign twf_m0_imag_val[511] = 9'sd98;

endmodule



